a0_0|NA|VAP
a0_0|NA|VAPs
a0_0|NA|vent acquired infection
a0_0|NA|vent acquired infections
a0_0|NA|vent acquired PNA
a0_0|NA|vent acquired PNAs
a0_0|NA|vent acquired pneumonias
a0_0|NA|vent acquired pneumonia
a0_0|NA|vent associated infection
a0_0|NA|vent associated infections
a0_0|NA|vent associated PNA
a0_0|NA|vent associated PNAs
a0_0|NA|vent associated pneumonia
a0_0|NA|vent associated pneumonias
a0_0|NA|vent infection
a0_0|NA|vent infections
a0_0|NA|vent PNA
a0_0|NA|vent PNAs
a0_0|NA|vent pneumonia
a0_0|NA|vent pneumonias
a0_0|NA|ventilator acquired infection
a0_0|NA|ventilator acquired infections
a0_0|NA|ventilator acquired PNA
a0_0|NA|ventilator acquired PNAs
a0_0|NA|ventilator acquired pneumonia
a0_0|NA|ventilator acquired pneumonias
a0_0|NA|ventilator associated infection
a0_0|NA|ventilator associated infections
a0_0|NA|ventilator infection
a0_0|NA|ventilator infections
a0_0|NA|ventilator PNA
a0_0|NA|ventilator PNAs
a0_0|NA|ventilator pneumonia
a0_0|NA|ventilator pneumonias
a0_0|NA|ventilator-associated PNA
a0_0|NA|ventilator-associated PNAs
a0_0|NA|ventilator-associated pneumonia
a0_0|NA|ventilator-associated pneumonias
a0_0|NA|ventilatory acquired infection
a0_0|NA|ventilatory acquired infections
a0_0|NA|ventilatory acquired PNA
a0_0|NA|ventilatory acquired PNAs
a0_0|NA|ventilatory acquired pneumonia
a0_0|NA|ventilatory acquired pneumonias
a0_0|NA|ventilatory associated infection
a0_0|NA|ventilatory infection
a0_0|NA|ventilatory infections
a0_0|NA|ventilatory PNA
a0_0|NA|ventilatory PNAs
a0_0|NA|ventilatory pneumonia
a0_0|NA|ventilatory pneumonias
a0_0|NA|ventilatory-associated PNA
a0_0|NA|ventilatory-associated PNAs
a0_0|NA|ventilatory-associated pneumonia
a0_0|NA|ventilatory-associated pneumonias
a0_0|NA|vent aquired pneumonia
a0_0|NA|ventilater-associated pneumonia
a0_1|NA|N95 respirator masks
a0_1|NA|N95 respirator mask
a0_1|NA|N95 respirators
a0_1|NA|N95 respirator
a0_1|NA|N95 masks
a0_1|NA|N95 mask
a0_1|NA|N95
a0_1|NA|N95s
a0_1|NA|N-95 respirator masks
a0_1|NA|N-95 respirator mask
a0_1|NA|N-95 respirators
a0_1|NA|N-95 respirator
a0_1|NA|N-95 masks
a0_1|NA|N-95 mask
a0_1|NA|N-95
a0_1|NA|N-95s
a0_2|NA|person-to-person transmission
a0_2|NA|human-to-human transmission
a0_2|NA|person-to-person transmissions
a0_2|NA|human-to-human transmissions
a0_2|NA|transmitted person-to-peson
a0_2|NA|transmitted human-to-human
a0_2|NA|transmitting person-to-peson
a0_2|NA|transmitting human-to-human
a0_2|NA|transmits person-to-peson
a0_2|NA|transmits human-to-human
a0_2|NA|transmit person-to-peson
a0_2|NA|transmit human-to-human
a0_2|NA|contagious disease
a0_2|NA|contagious diseases
a0_2|NA|contagiousness
a0_2|NA|contagious
a0_3|NA|first human drug trial
a0_3|NA|first human drug trials
a0_3|NA|human drug trial
a0_3|NA|human drug trials
a0_3|NA|first drug trial in humans
a0_3|NA|first drug trials in humans
a0_3|NA|drug trial in humans
a0_3|NA|drug trials in humans
a0_3|NA|drug trial
a0_3|NA|drug trials
a0_4|NA|U07.1
a0_4|NA|COVID-19
a0_4|NA|COVID19
a0_5|NA|vaccine design
a0_5|NA|vaccine designs
a0_5|NA|vaccine research
a0_5|NA|design of vaccines
a0_5|NA|design of vaccination
a0_5|NA|designing vaccines
a0_5|NA|designed vaccines
a0_5|NA|designs vaccines
a0_5|NA|design vaccines
a0_5|NA|designing the vaccine
a0_5|NA|designed the vaccine
a0_5|NA|designs the vaccine
a0_5|NA|design the vaccine
a0_5|NA|designing a vaccine
a0_5|NA|designed a vaccine
a0_5|NA|designs a vaccine
a0_5|NA|design a vaccine
a0_6|NA|COVID-19 Ab IgM
a0_6|NA|COVID-19 Ab immunoglobulin M
a0_6|NA|COVID-19 antibody IgM
a0_6|NA|COVID-19 antibody immunoglobulin M
a0_6|NA|COVID-19 Ab
a0_6|NA|COVID-19 Abs
a0_6|NA|COVID-19 antibodies
a0_6|NA|COVID-19 antibody
a0_6|NA|immunoglobulin M COVID-19
a0_6|NA|IgM COVID-19
a0_6|NA|immunoglobulin M to COVID-19
a0_6|NA|IgM to COVID-19
a0_6|NA|antibodies to COVID-19
a0_6|NA|antibody to COVID-19
a0_6|NA|Abs to COVID-19
a0_6|NA|Ab to COVID-19
a0_6|NA|COVID19 Ab IgM
a0_6|NA|COVID19 Ab immunoglobulin M
a0_6|NA|COVID19 antibody IgM
a0_6|NA|COVID19 antibody immunoglobulin M
a0_6|NA|COVID19 Ab
a0_6|NA|COVID19 Abs
a0_6|NA|COVID19 antibodies
a0_6|NA|COVID19 antibody
a0_6|NA|immunoglobulin M COVID19
a0_6|NA|IgM COVID19
a0_6|NA|immunoglobulin M to COVID19
a0_6|NA|IgM to COVID19
a0_6|NA|antibodies to COVID19
a0_6|NA|antibody to COVID19
a0_6|NA|Abs to COVID19
a0_6|NA|Ab to COVID19
a0_6|NA|COVID Ab IgM
a0_6|NA|COVID Ab immunoglobulin M
a0_6|NA|COVID antibody IgM
a0_6|NA|COVID antibody immunoglobulin M
a0_6|NA|COVID Ab
a0_6|NA|COVID Abs
a0_6|NA|COVID antibodies
a0_6|NA|COVID antibody
a0_6|NA|immunoglobulin M COVID
a0_6|NA|IgM COVID
a0_6|NA|immunoglobulin M to COVID
a0_6|NA|IgM to COVID
a0_6|NA|antibodies to COVID
a0_6|NA|antibody to COVID
a0_6|NA|Abs to COVID
a0_6|NA|Ab to COVID
a0_6|NA|coronavirus Ab IgM
a0_6|NA|coronavirus Ab immunoglobulin M
a0_6|NA|coronavirus antibody IgM
a0_6|NA|coronavirus antibody immunoglobulin M
a0_6|NA|coronavirus Ab
a0_6|NA|coronavirus Abs
a0_6|NA|coronavirus antibodies
a0_6|NA|coronavirus antibody
a0_6|NA|immunoglobulin M coronavirus
a0_6|NA|IgM coronavirus
a0_6|NA|immunoglobulin M to coronavirus
a0_6|NA|IgM to coronavirus
a0_6|NA|antibodies to coronavirus
a0_6|NA|antibody to coronavirus
a0_6|NA|Abs to coronavirus
a0_6|NA|Ab to coronavirus
a0_6|NA|immunoglobulin M to the coronavirus
a0_6|NA|IgM to the coronavirus
a0_6|NA|antibodies to the coronavirus
a0_6|NA|antibody to the coronavirus
a0_6|NA|Abs to the coronavirus
a0_6|NA|Ab to the coronavirus
a0_6|NA|immunoglobulin M to the novel coronavirus
a0_6|NA|IgM to the novel coronavirus
a0_6|NA|antibodies to the novel coronavirus
a0_6|NA|antibody to the novel coronavirus
a0_6|NA|Abs to the novel coronavirus
a0_6|NA|Ab to the novel coronavirus
a0_7|NA|N95 respirator masks
a0_7|NA|N95 respirator mask
a0_7|NA|N95 respirators
a0_7|NA|N95 respirator
a0_7|NA|N95 masks
a0_7|NA|N95 mask
a0_7|NA|respirator masks
a0_7|NA|respirator mask
a0_8|NA|COVID-19 death toll
a0_8|NA|COVID-19 death tolls
a0_8|NA|COVID-19 mortality
a0_8|NA|COVID-19 deaths
a0_8|NA|COVID-19 death
a0_8|NA|COVID19 deaths
a0_8|NA|COVID19 death
a0_8|NA|COVID deaths
a0_8|NA|COVID death
a0_8|NA|coronavirus-19 deaths
a0_8|NA|coronavirus-19 death
a0_8|NA|deaths from COVID-19
a0_8|NA|death from COVID-19
a0_8|NA|dying from COVID-19
a0_8|NA|died from COVID-19
a0_8|NA|COVID19 death toll
a0_8|NA|COVID19 death tolls
a0_8|NA|COVID19 mortality
a0_8|NA|deaths from COVID19
a0_8|NA|death from COVID19
a0_8|NA|dying from COVID19
a0_8|NA|died from COVID19
a0_8|NA|COVID death toll
a0_8|NA|COVID death tolls
a0_8|NA|COVID mortality
a0_8|NA|deaths from COVID
a0_8|NA|death from COVID
a0_8|NA|dying from COVID
a0_8|NA|died from COVID
a0_8|NA|coronavirus death toll
a0_8|NA|coronavirus death tolls
a0_8|NA|coronavirus mortality
a0_8|NA|deaths from coronavirus
a0_8|NA|death from coronavirus
a0_8|NA|dying from coronavirus
a0_8|NA|died from coronavirus
a0_9|NA|COVID-19 symptom
a0_9|NA|COVID-19 symptoms
a0_9|NA|symptom of COVID-19
a0_9|NA|symptoms of COVID-19
a0_9|NA|symptomatic COVID-19
a0_9|NA|COVID19 symptom
a0_9|NA|COVID19 symptoms
a0_9|NA|symptom of COVID19
a0_9|NA|symptoms of COVID19
a0_9|NA|symptomatic COVID19
a0_9|NA|COVID symptom
a0_9|NA|COVID symptoms
a0_9|NA|symptom of COVID
a0_9|NA|symptoms of COVID
a0_9|NA|symptomatic COVID
a0_9|NA|coronavirus symptom
a0_9|NA|coronavirus symptoms
a0_9|NA|symptom of coronavirus
a0_9|NA|symptoms of coronavirus
a0_9|NA|symptomatic coronavirus
a0_11|NA|KN95 masks
a0_11|NA|KN95 mask
a0_11|NA|N95 masks
a0_11|NA|N95 mask
a0_11|NA|KN-95 masks
a0_11|NA|KN-95 mask
a0_11|NA|N-95 masks
a0_11|NA|N-95 mask
a0_11|NA|KN95 protection mask
a0_11|NA|KN95 protection masks
a0_11|NA|KN95
a0_11|NA|N95
a0_12|NA|paediatric inflammatory multisystem syndrome
a0_12|NA|pediatric inflammatory multisystem syndrome
a0_12|NA|paediatric inflammatory multi-system syndrome
a0_12|NA|pediatric inflammatory multi-system syndrome
a0_12|NA|pediatric inflammatory myocardial syndrome
a0_12|NA|paediatric inflammatory myocardial syndrome
a0_12|NA|PIMS
a0_12|NA|PIMS-TS
a0_13|NA|ventilator-dependent pneumonia
a0_13|NA|ventilator associated pneumonia
a0_13|NA|ventilator-dependent PNA
a0_13|NA|ventilator associated PNA
a0_13|NA|ventilator-dependent
a0_13|NA|ventilater-dependent pneumonia
a0_13|NA|ventilater associated pneumonia
a0_13|NA|ventilater-dependent PNA
a0_13|NA|ventilater associated PNA
a0_13|NA|pneumonia
a0_14|NA|hydroxychloroquine
a0_14|NA|Plaquenil sulfate
a0_14|NA|Plaquenil
a0_14|NA|anti-malarial
a0_15|NA|chloroquine
a0_15|NA|Aralen
a0_15|NA|anti-malarial
a0_15|NA|chlororquine
a0_15|NA|choroquine
a0_15|NA|hloroquine
a0_15|NA|chloroqunie
a0_15|NA|chloraquine
a0_15|NA|choloroquine
a0_15|NA|ochloroquine
a0_15|NA|chlroroquine
a0_15|NA|chlroquine
a0_15|NA|chlorquine
a0_15|NA|cholroquine
a0_15|NA|chloroquin
a0_15|NA|chloroquines
a0_15|NA|chloroqine
a0_15|NA|chloroxuine
a0_15|NA|chloriquine
a0_15|NA|chloroguine
a0_15|NA|chloroquinie
a0_15|NA|cloroquine
a0_15|NA|chrloroquine
a0_16|NA|Pediatric Inflammatory Myocardial Syndrome
a0_16|NA|Kawasaki-like condition
a0_16|NA|Kawasaki-like syndrome
a0_16|NA|Kawasaki-like illness
a0_16|NA|COVID-related Kawasaki like illness
a0_16|NA|COVID-related Kawasaki like syndrome
a0_16|NA|COVID-related Kawasaki like disease
a0_16|NA|COVID19-related Kawasaki like illness
a0_16|NA|COVID19-related Kawasaki like syndrome
a0_16|NA|COVID10-related Kawasaki like disease
a0_16|NA|COVID-19-related Kawasaki like illness
a0_16|NA|COVID-19-related Kawasaki like syndrome
a0_16|NA|COVID-19-related Kawasaki like disease
a0_16|NA|coronavirus-related Kawasaki like illness
a0_16|NA|coronavirus-related Kawasaki like syndrome
a0_16|NA|coronavirus-related Kawasaki like disease
a0_16|NA|Pediatric Inflammatory Myocardial Syndromes
a0_16|NA|Kawasaki-like conditions
a0_16|NA|Kawasaki-like syndromes
a0_16|NA|Kawasaki-like illnesses
a0_16|NA|COVID-related Kawasaki like illnesses
a0_16|NA|COVID-related Kawasaki like syndromes
a0_16|NA|COVID-related Kawasaki like diseases
a0_16|NA|COVID19-related Kawasaki like illnesses
a0_16|NA|COVID19-related Kawasaki like syndromes
a0_16|NA|COVID10-related Kawasaki like diseases
a0_16|NA|COVID-19-related Kawasaki like illnesses
a0_16|NA|COVID-19-related Kawasaki like syndromes
a0_16|NA|COVID-19-related Kawasaki like diseases
a0_16|NA|coronavirus-related Kawasaki like illnesses
a0_16|NA|coronavirus-related Kawasaki like syndromes
a0_16|NA|coronavirus-related Kawasaki like diseases
a0_16|NA|Kawasaki disease-like condition
a0_16|NA|Kawasaki disease-like syndrome
a0_16|NA|Kawasaki disease-like illness
a0_16|NA|COVID-related Kawasaki disease like illness
a0_16|NA|COVID-related Kawasaki disease like syndrome
a0_16|NA|COVID19-related Kawasaki disease like illness
a0_16|NA|COVID19-related Kawasaki disease like syndrome
a0_16|NA|COVID-19-related Kawasaki disease like illness
a0_16|NA|COVID-19-related Kawasaki disease like syndrome
a0_16|NA|coronavirus-related Kawasaki disease like illness
a0_16|NA|coronavirus-related Kawasaki disease like syndromeKawasaki disease-like conditions
a0_16|NA|Kawasaki disease-like syndromes
a0_16|NA|Kawasaki disease-like illnesses
a0_16|NA|COVID-related Kawasaki disease like illnesses
a0_16|NA|COVID-related Kawasaki disease like syndromes
a0_16|NA|COVID19-related Kawasaki disease like illnesses
a0_16|NA|COVID19-related Kawasaki disease like syndromes
a0_16|NA|COVID-19-related Kawasaki disease like illnesses
a0_16|NA|COVID-19-related Kawasaki disease like syndromes
a0_16|NA|coronavirus-related Kawasaki disease like illnesses
a0_16|NA|coronavirus-related Kawasaki disease like syndromes
a0_17|NA|nasopharyngeal swabs
a0_17|NA|nasopharyngeal swab
a0_17|NA|nasopharyngeal sample
a0_17|NA|nasopharyngeal samples
a0_17|NA|nasopharyngeal sampling
a0_17|NA|naso-pharyngeal swabs
a0_17|NA|naso-pharyngeal swab
a0_17|NA|naso-pharyngeal sample
a0_17|NA|naso-pharyngeal samples
a0_17|NA|naso-pharyngeal sampling
a0_17|NA|nasopharynx swabs
a0_17|NA|nasopharynx swab
a0_17|NA|nasopharynx sample
a0_17|NA|nasopharynx samples
a0_17|NA|nasopharynx sampling
a0_17|NA|naso-pharynx swabs
a0_17|NA|naso-pharynx swab
a0_17|NA|naso-pharynx sample
a0_17|NA|naso-pharynx samples
a0_17|NA|naso-pharynx sampling
a0_17|NA|NP swabs
a0_17|NA|NP swab
a0_17|NA|NP sample
a0_17|NA|NP samples
a0_17|NA|NP sampling
a0_17|NA|swabbing the NP
a0_17|NA|swabbing the naso-pharynx
a0_17|NA|swabbing the nasopharynx
a0_17|NA|swabbed the NP
a0_17|NA|swabbed the naso-pharynx
a0_17|NA|swabbed the nasopharynx
a0_17|NA|swabs the NP
a0_17|NA|swabs the naso-pharynx
a0_17|NA|swabs the nasopharynx
a0_17|NA|swab the NP
a0_17|NA|swab the naso-pharynx
a0_17|NA|swab the nasopharynx
a0_17|NA|samples from the NP
a0_17|NA|sample from the NP
a0_17|NA|samples from NP
a0_17|NA|sample from NP
a0_17|NA|samples from the nasopharynx
a0_17|NA|sample from the nasopharynx
a0_17|NA|samples from nasopharynx
a0_17|NA|sample from nasopharynx
a0_17|NA|samples from the naso-pharynx
a0_17|NA|sample from the naso-pharynx
a0_17|NA|samples from naso-pharynx
a0_17|NA|sample from naso-pharynx
a0_17|NA|sampling the NP
a0_17|NA|sampled the NP
a0_17|NA|samples the NP
a0_17|NA|sample the NP
a0_17|NA|sampling the nasopharynx
a0_17|NA|sampled the nasopharynx
a0_17|NA|samples the nasopharynx
a0_17|NA|sample the nasopharynx
a0_17|NA|sampling the naso-pharynx
a0_17|NA|sampled the naso-pharynx
a0_17|NA|samples the naso-pharynx
a0_17|NA|sample the naso-pharynx
a0_18|NA|COVID-19 antibodies
a0_18|NA|COVID-19 Abs
a0_18|NA|COVID-19 antibody
a0_18|NA|COVID-19 antibody testing
a0_18|NA|COVID-19 antibody tests
a0_18|NA|COVID-19 antibody test
a0_18|NA|COVID-19 Ab
a0_18|NA|COVID-19 Ab testing
a0_18|NA|COVID-19 Ab tests
a0_18|NA|COVID-19 Ab test
a0_18|NA|COVID19 antibodies
a0_18|NA|COVID19 Abs
a0_18|NA|COVID19 antibody
a0_18|NA|COVID19 antibody testing
a0_18|NA|COVID19 antibody tests
a0_18|NA|COVID19 antibody test
a0_18|NA|COVID19 Ab
a0_18|NA|COVID19 Ab testing
a0_18|NA|COVID19 Ab tests
a0_18|NA|COVID19 Ab test
a0_18|NA|COVID antibodies
a0_18|NA|COVID Abs
a0_18|NA|COVID antibody
a0_18|NA|COVID antibody testing
a0_18|NA|COVID antibody tests
a0_18|NA|COVID antibody test
a0_18|NA|COVID Ab
a0_18|NA|COVID Ab testing
a0_18|NA|COVID Ab tests
a0_18|NA|COVID Ab test
a0_18|NA|testing for COVID-19 antibodies
a0_18|NA|testing for COVID-19 Abs
a0_18|NA|testing for COVID-19 antibody
a0_18|NA|testing for COVID-19 Ab
a0_18|NA|tested for COVID-19 antibodies
a0_18|NA|tested for COVID-19 Abs
a0_18|NA|tested for COVID-19 antibody
a0_18|NA|tested for COVID-19 Ab
a0_18|NA|tests for COVID-19 antibodies
a0_18|NA|tests for COVID-19 Abs
a0_18|NA|tests for COVID-19 antibody
a0_18|NA|tests for COVID-19 Ab
a0_18|NA|test for COVID-19 antibodies
a0_18|NA|test for COVID-19 Abs
a0_18|NA|test for COVID-19 antibody
a0_18|NA|test for COVID-19 Ab
a0_18|NA|testing for COVID19 antibodies
a0_18|NA|testing for COVID19 Abs
a0_18|NA|testing for COVID19 antibody
a0_18|NA|testing for COVID19 Ab
a0_18|NA|tested for COVID19 antibodies
a0_18|NA|tested for COVID19 Abs
a0_18|NA|tested for COVID19 antibody
a0_18|NA|tested for COVID19 Ab
a0_18|NA|tests for COVID19 antibodies
a0_18|NA|tests for COVID19 Abs
a0_18|NA|tests for COVID19 antibody
a0_18|NA|tests for COVID19 Ab
a0_18|NA|test for COVID19 antibodies
a0_18|NA|test for COVID19 Abs
a0_18|NA|test for COVID19 antibody
a0_18|NA|test for COVID19 Ab
a0_18|NA|testing for COVID antibodies
a0_18|NA|testing for COVID Abs
a0_18|NA|testing for COVID antibody
a0_18|NA|testing for COVID Ab
a0_18|NA|tested for COVID antibodies
a0_18|NA|tested for COVID Abs
a0_18|NA|tested for COVID antibody
a0_18|NA|tested for COVID Ab
a0_18|NA|tests for COVID antibodies
a0_18|NA|tests for COVID Abs
a0_18|NA|tests for COVID antibody
a0_18|NA|tests for COVID Ab
a0_18|NA|test for COVID antibodies
a0_18|NA|test for COVID Abs
a0_18|NA|test for COVID antibody
a0_18|NA|test for COVID Ab
a0_18|NA|COVID-19
a0_18|NA|COVID19
a0_19|NA|Pediatric Inflammatory Myocardial Syndrome
a0_19|NA|COVID-19
a0_20|NA|COVID-19 case
a0_20|NA|COVID19 case
a0_20|NA|COVID case
a0_20|NA|coronavirus case
a0_20|NA|COVID-19 diagnosis
a0_20|NA|COVID19 diagnosis
a0_20|NA|COVID diagnosis
a0_20|NA|coronavirus diagnosis
a0_20|NA|positive for COVID-19
a0_20|NA|positive for COVID19
a0_20|NA|positive for COVID
a0_20|NA|positive for coronavirus
a0_20|NA|positive COVID-19
a0_20|NA|positive COVID19
a0_20|NA|positive COVID
a0_20|NA|positive coronavirus
a0_21|NA|Plaquenil
a0_21|NA|plaquinal
a0_21|NA|plaquneil
a0_21|NA|placquenil
a0_21|NA|plaqyenil
a0_21|NA|plaqueuil
a0_21|NA|plaqueniil
a0_21|NA|plaqunenil
a0_21|NA|plaqucnil
a0_21|NA|plaqueneil
a0_21|NA|plaquemil
a0_21|NA|plaquenail
a0_21|NA|plaqueenil
a0_21|NA|plaguenil
a0_21|NA|plaquenol
a0_21|NA|plazuenil
a0_21|NA|plaquenily
a0_21|NA|plaqueinil
a0_21|NA|plauquenil
a0_21|NA|plaquenil1
a0_21|NA|dplaquenil
a0_21|NA|dlaquenil
a0_21|NA|pplaquenil
a0_21|NA|plaqueninl
a0_21|NA|plaqenil
a0_21|NA|planquenil
a0_21|NA|plaquonil
a0_21|NA|plaqunil
a0_21|NA|oplaquenil
a0_21|NA|plaqueinl
a0_21|NA|plquenil
a0_21|NA|plaqqenil
a0_21|NA|plaqquenil
a0_21|NA|plaquenuil
a0_21|NA|plaquelnil
a0_21|NA|plagquenil
a0_21|NA|plaquenial
a0_21|NA|plaqienil
a0_21|NA|plaquenal
a0_21|NA|plqauenil
a0_21|NA|plaquennil
a0_21|NA|plaquenel
a0_21|NA|plaqueil
a0_21|NA|plaqueril
a0_21|NA|plaquanil
a0_21|NA|laquenil
a0_21|NA|plaequenil
a0_21|NA|plaqusenil
a0_21|NA|plaquenfil
a0_21|NA|plaquenbil
a0_21|NA|plaquenic
a0_21|NA|plawuenil
a0_21|NA|cplaquenil
a0_21|NA|paquenil
a0_21|NA|plaquenul
a0_21|NA|plaquenyl
a0_21|NA|palquenil
a0_21|NA|plaquienil
a0_21|NA|plequenil
a0_21|NA|plaquenils
a0_21|NA|plaquenl
a0_21|NA|plaquenilt
a0_21|NA|plqquenil
a0_21|NA|plaqueunil
a0_21|NA|plaquenili
a0_21|NA|praquenil
a0_21|NA|plaquenilk
a0_21|NA|plaquenill
a0_21|NA|plaquenile
a0_21|NA|plasquenil
a0_21|NA|plaqueni
a0_21|NA|plaqeunil
a0_21|NA|plaquinil
a0_21|NA|plalquenil
a0_21|NA|plaquenitl
a0_21|NA|plaqnenil
a0_21|NA|plauqenil
a0_21|NA|plauenil
a0_21|NA|plaquentil
a0_21|NA|plaqvenil
a0_21|NA|plaquenicl
a0_21|NA|plaquenix
a0_21|NA|plaquenril
a0_22|NA|social distancing
a0_22|NA|social distance
a0_22|NA|social distancers
a0_22|NA|social distancer
a0_22|NA|socially distancing
a0_22|NA|socially distanced
a0_22|NA|socially distances
a0_22|NA|socially distance
a0_22|NA|6 feet apart
a0_22|NA|6 feet away
a0_22|NA|fix feet apart
a0_22|NA|six feet away
a0_22|NA|2 meters apart
a0_22|NA|2 meters away
a0_22|NA|two meters apart
a0_22|NA|two meters away
a0_22|NA|socialdistancing
a0_23|NA|COVID-19 pandemic
a0_23|NA|COVID19 pandemic
a0_23|NA|COVID pandemic
a0_23|NA|coronavirus pandemic
a0_23|NA|COVID-19 crisis
a0_23|NA|COVID19 crisis
a0_23|NA|COVID crisis
a0_23|NA|coronavirus crisis
a0_23|NA|COVID-19 crises
a0_23|NA|COVID19 crises
a0_23|NA|COVID crises
a0_23|NA|coronavirus crises
a0_23|NA|COVID-19 situation
a0_23|NA|COVID19 situation
a0_23|NA|COVID situation
a0_23|NA|coronavirus situation
a0_23|NA|COVID-19 situations
a0_23|NA|COVID19 situations
a0_23|NA|COVID situations
a0_23|NA|coronavirus situations
a0_24|NA|contact tracing
a0_24|NA|tracing her contacts
a0_24|NA|tracing his contacts
a0_24|NA|tracing the contacts
a0_24|NA|tracing contacts
a0_24|NA|close contact tracing
a0_24|NA|tracing her close contacts
a0_24|NA|tracing his close contacts
a0_24|NA|tracing the close contacts
a0_24|NA|tracing close contacts
a0_24|NA|traced her contacts
a0_24|NA|traced his contacts
a0_24|NA|traced the contacts
a0_24|NA|traced contacts
a0_24|NA|traced her close contacts
a0_24|NA|traced his close contacts
a0_24|NA|traced the close contacts
a0_24|NA|traced close contacts
a0_24|NA|traces her contacts
a0_24|NA|traces his contacts
a0_24|NA|traces the contacts
a0_24|NA|traces contacts
a0_24|NA|traces her close contacts
a0_24|NA|traces his close contacts
a0_24|NA|traces the close contacts
a0_24|NA|traces close contacts
a0_24|NA|trace her contacts
a0_24|NA|trace his contacts
a0_24|NA|trace the contacts
a0_24|NA|trace contacts
a0_24|NA|trace her close contacts
a0_24|NA|trace his close contacts
a0_24|NA|trace the close contacts
a0_24|NA|trace close contacts
a0_25|NA|artificial respiration
a0_25|NA|artificial respirators
a0_25|NA|artificial respirator
a0_25|NA|artificial ventilation
a0_25|NA|artificial ventilators
a0_25|NA|artificial ventilator
a0_25|NA|artificially ventilating
a0_25|NA|artificially ventilated
a0_25|NA|artificially ventilates
a0_25|NA|artificially ventilate
a0_25|NA|breathing machines
a0_25|NA|breathing machine
a0_25|NA|mechanically ventilated
a0_25|NA|mechanical ventilation
a0_25|NA|mechanical ventilators
a0_25|NA|mechanical ventilator
a0_25|NA|mechanical vents
a0_25|NA|mechanical vent
a0_25|NA|ventilations
a0_25|NA|ventilation
a0_25|NA|ventilators
a0_25|NA|ventilator
a0_25|NA|ventilating
a0_25|NA|ventilated
a0_25|NA|ventilates
a0_25|NA|ventilate
a0_25|NA|vented
a0_25|NA|on a ventilator
a0_25|NA|on a vent
a0_25|NA|on ventilator
a0_25|NA|on vent
a0_25|NA|vents
a0_25|NA|vent
a0_25|NA|ventilatin
a0_25|NA|ventillation
a0_25|NA|ventailation
a0_25|NA|ventialltion
a0_25|NA|ventalation
a0_25|NA|ventliation
a0_25|NA|ventilater
a0_25|NA|ventalator
a0_25|NA|ventelator
a0_25|NA|ventillator
a0_25|NA|ventalotor
a0_25|NA|ventialtion
a0_25|NA|venntilat
a0_25|NA|ventilato
a0_25|NA|ventilatory
a0_25|NA|venilation
a0_25|NA|ventilaiton
a0_25|NA|ventilaor
a0_25|NA|ventilatio
a0_25|NA|ventilatioin
a0_25|NA|ventilat
a0_25|NA|vetilator
a0_25|NA|mechanical ventillation
a0_25|NA|mechnical ventilation
a0_25|NA|ventilaton
a0_25|NA|ventialtor
a0_25|NA|ventilacion
a0_25|NA|ventilantion
a0_25|NA|ventalated
a0_25|NA|ventilarot
a0_25|NA|ventilationa
a0_25|NA|venitlator
a0_25|NA|ventilaotr
a0_25|NA|ventilatro
a0_25|NA|ventiltaor
a0_25|NA|ventliator
a0_25|NA|vnetilator
a0_25|NA|veantilator
a0_25|NA|veintilator
a0_25|NA|venatilator
a0_25|NA|venetilator
a0_25|NA|venitilator
a0_25|NA|ventailator
a0_25|NA|ventiilator
a0_25|NA|ventilaator
a0_25|NA|ventilaotor
a0_25|NA|ventilataor
a0_25|NA|ventilateor
a0_25|NA|ventilatior
a0_25|NA|ventilatoar
a0_25|NA|ventilatoer
a0_25|NA|ventilatoir
a0_25|NA|ventilatoor
a0_25|NA|ventilatore
a0_25|NA|ventilatorr
a0_25|NA|ventilatoru
a0_25|NA|ventilatr
a0_25|NA|ventilattor
a0_25|NA|ventiliator
a0_25|NA|ventiloator
a0_25|NA|ventiltor
a0_25|NA|ventiolator
a0_25|NA|ventiulator
a0_25|NA|ventlator
a0_25|NA|venttilator
a0_25|NA|ventuilator
a0_25|NA|ventyilator
a0_25|NA|vewntilator
a0_25|NA|vntilator
a0_25|NA|vventilator
a0_25|NA|vwentilator
a0_25|NA|fentilator
a0_25|NA|vantilator
a0_25|NA|ventilador
a0_25|NA|ventilatir
a0_25|NA|ventilitor
a0_25|NA|ventilltor
a0_25|NA|ventilotor
a0_25|NA|ventllator
a0_25|NA|ventolator
a0_25|NA|ventulator
a0_25|NA|evntilator
a0_25|NA|vetnilator
a0_25|NA|ventiator
a0_25|NA|nventilator
a0_25|NA|ventiltator
a0_25|NA|venthilator
a0_25|NA|ventialator
a0_25|NA|ventilartor
a0_25|NA|entilator
a0_25|NA|verntilator
a0_25|NA|ventilaltor
a0_25|NA|ventlilator
a0_25|NA|ventilatlor
a0_25|NA|rventilator
a0_25|NA|ventinlator
a0_25|NA|venilator
a0_25|NA|ventilatord
a0_25|NA|ventilatort
a0_25|NA|aventilator
a0_25|NA|eventilator
a0_25|NA|oventilator
a0_25|NA|ventilatorl
a0_25|NA|vlentilator
a0_25|NA|ventrilator
a0_25|NA|ventilatorx
a0_25|NA|ventitlator
a0_25|NA|vetntilator
a0_25|NA|vemntilator
a0_25|NA|pventilator
a0_25|NA|ventilatot
a0_25|NA|ventilatos
a0_25|NA|ventilztor
a0_25|NA|vemtilator
a0_25|NA|wentilator
a0_25|NA|vertilator
a0_25|NA|hentilator
a0_25|NA|ventilaror
a0_25|NA|ventilatoe
a0_25|NA|ventilatoy
a0_25|NA|bentilator
a0_25|NA|ventrlator
a0_25|NA|veitilator
a0_25|NA|vebtilator
a0_25|NA|ventilatpr
a0_25|NA|ventitator
a0_25|NA|ventirator
a0_25|NA|centilator
a0_25|NA|venrilator
a0_25|NA|venitlation
a0_25|NA|vnetilation
a0_25|NA|veentilation
a0_25|NA|venatilation
a0_25|NA|venetilation
a0_25|NA|venitilation
a0_25|NA|venntilation
a0_25|NA|ventiilation
a0_25|NA|ventilaation
a0_25|NA|ventilaition
a0_25|NA|ventilation1
a0_25|NA|ventilationi
a0_25|NA|ventilationo
a0_25|NA|ventilationw
a0_25|NA|ventiliation
a0_25|NA|ventiltion
a0_25|NA|ventiolation
a0_25|NA|ventiulation
a0_25|NA|ventlation
a0_25|NA|venttilation
a0_25|NA|ventuilation
a0_25|NA|vntilation
a0_25|NA|vventilation
a0_25|NA|fentilation
a0_25|NA|vantilation
a0_25|NA|ventelation
a0_25|NA|ventilition
a0_25|NA|ventllation
a0_25|NA|ventolation
a0_25|NA|ventulation
a0_25|NA|ventilatino
a0_25|NA|ventilatoin
a0_25|NA|ventiltaion
a0_25|NA|ventiation
a0_25|NA|venticlation
a0_25|NA|ventiklation
a0_25|NA|ventilaion
a0_25|NA|venbtilation
a0_25|NA|ventialation
a0_25|NA|ventiltation
a0_25|NA|vbentilation
a0_25|NA|ventilartion
a0_25|NA|vdentilation
a0_25|NA|velntilation
a0_25|NA|ventilaltion
a0_25|NA|ventlilation
a0_25|NA|ventilatgion
a0_25|NA|rventilation
a0_25|NA|vetilation
a0_25|NA|vemntilation
a0_25|NA|mventilation
a0_25|NA|venrtilation
a0_25|NA|ventrilation
a0_25|NA|ventilataion
a0_25|NA|ventilatiion
a0_25|NA|ventilatiojn
a0_25|NA|ventilatioon
a0_25|NA|ventilatiuon
a0_25|NA|ventilatoion
a0_25|NA|ventilattion
a0_25|NA|ventilatuion
a0_25|NA|ventilatyion
a0_25|NA|ventilatrion
a0_25|NA|ventinlation
a0_25|NA|ventilastion
a0_25|NA|ventilaztion
a0_25|NA|vevntilation
a0_25|NA|verntilation
a0_25|NA|vrentilation
a0_25|NA|aventilation
a0_25|NA|eventilation
a0_25|NA|oventilation
a0_25|NA|ventilationz
a0_25|NA|ventilationm
a0_25|NA|ventilationl
a0_25|NA|ventilationg
a0_25|NA|venmtilation
a0_25|NA|vcentilation
a0_25|NA|ventitlation
a0_25|NA|entilation
a0_25|NA|mentilation
a0_25|NA|ventilaaion
a0_25|NA|vertilation
a0_25|NA|ventitation
a0_25|NA|vdntilation
a0_25|NA|gentilation
a0_25|NA|centilation
a0_25|NA|vemtilation
a0_25|NA|ventilatiom
a0_25|NA|ventilasion
a0_25|NA|ventilstion
a0_25|NA|ventilarion
a0_25|NA|ventication
a0_25|NA|wentilation
a0_25|NA|venitlated
a0_25|NA|ventiltaed
a0_25|NA|ventliated
a0_25|NA|vnetilated
a0_25|NA|venitilated
a0_25|NA|ventailated
a0_25|NA|ventiilated
a0_25|NA|ventilataed
a0_25|NA|ventilatedt
a0_25|NA|ventilatied
a0_25|NA|ventilatoed
a0_25|NA|ventilhated
a0_25|NA|ventiliated
a0_25|NA|ventillated
a0_25|NA|ventilted
a0_25|NA|ventlated
a0_25|NA|venttilated
a0_25|NA|vewntilated
a0_25|NA|fentilated
a0_25|NA|vantilated
a0_25|NA|ventelated
a0_25|NA|ventillted
a0_25|NA|ventolated
a0_25|NA|ventulated
a0_25|NA|ventialted
a0_25|NA|vetnilated
a0_25|NA|ventiated
a0_25|NA|ventiltated
a0_25|NA|ventilateds
a0_25|NA|ventilatedl
a0_25|NA|ventialated
a0_25|NA|entilated
a0_25|NA|vrentilated
a0_25|NA|rventilated
a0_25|NA|venilated
a0_25|NA|eventilated
a0_25|NA|oventilated
a0_25|NA|ventilaed
a0_25|NA|ventilatd
a0_25|NA|ventrilated
a0_25|NA|ventitlated
a0_25|NA|vetilated
a0_25|NA|venmtilated
a0_25|NA|ventilatec
a0_25|NA|vestilated
a0_25|NA|vemtilated
a0_25|NA|vertilated
a0_25|NA|ventilared
a0_25|NA|vnt
a0_25|NA|vnet
a0_26|NA|COVID 19 test result presumed positive
a0_26|NA|COVID19 test result presumed positive
a0_26|NA|COVID 19 test presumed positive
a0_26|NA|COVID19 test presumed positive
a0_26|NA|COVID 19 presumed positive
a0_26|NA|COVID19 presumed positive
a0_26|NA|presumptive positive COVID 19 test result
a0_26|NA|presumptive positive COVID 19 result
a0_26|NA|presumptive positive COVID19 test result
a0_26|NA|presumptive positive COVID19 result
a0_26|NA|presumptive positive COVID test result
a0_26|NA|presumptive positive COVID result
a0_26|NA|presumptive positive for 2019 novel coronavirus
a0_26|NA|presumptive positive for novel coronavirus
a0_26|NA|presumptive positive for COVID 19
a0_26|NA|presumptive positive for COVID19
a0_26|NA|presumptive positive for COVID
a0_26|NA|presumptive positive for 2019 novel coronavirus RNA
a0_26|NA|presumptive positive for novel coronavirus RNA
a0_26|NA|presumptive positive for COVID 19 RNA
a0_26|NA|presumptive positive for COVID19 RNA
a0_26|NA|COVID 19 test result presumed pos
a0_26|NA|COVID19 test result presumed pos
a0_26|NA|COVID 19 test presumed pos
a0_26|NA|COVID19 test presumed pos
a0_26|NA|COVID 19 presumed pos
a0_26|NA|COVID19 presumed pos
a0_26|NA|presumptive pos COVID 19 test result
a0_26|NA|presumptive pos COVID 19 result
a0_26|NA|presumptive pos COVID19 test result
a0_26|NA|presumptive pos COVID19 result
a0_26|NA|presumptive pos COVID test result
a0_26|NA|presumptive pos COVID result
a0_26|NA|presumptive pos for 2019 novel coronavirus
a0_26|NA|presumptive pos for novel coronavirus
a0_26|NA|presumptive pos for COVID 19
a0_26|NA|presumptive pos for COVID19
a0_26|NA|presumptive pos for COVID
a0_26|NA|presumptive pos for 2019 novel coronavirus RNA
a0_26|NA|presumptive pos for novel coronavirus RNA
a0_26|NA|presumptive pos for COVID 19 RNA
a0_26|NA|presumptive pos for COVID19 RNA
a0_26|NA|presumed positive COVID 19 test result
a0_26|NA|presumed positive COVID 19 result
a0_26|NA|presumed positive COVID19 test result
a0_26|NA|presumed positive COVID19 result
a0_26|NA|presumed positive COVID test result
a0_26|NA|presumed positive COVID result
a0_26|NA|presumed positive for 2019 novel coronavirus
a0_26|NA|presumed positive for novel coronavirus
a0_26|NA|presumed positive for COVID 19
a0_26|NA|presumed positive for COVID19
a0_26|NA|presumed positive for COVID
a0_26|NA|presumed positive for 2019 novel coronavirus RNA
a0_26|NA|presumed positive for novel coronavirus RNA
a0_26|NA|presumed positive for COVID 19 RNA
a0_26|NA|presumed positive for COVID19 RNA
a0_26|NA|presumed pos COVID 19 test result
a0_26|NA|presumed pos COVID 19 result
a0_26|NA|presumed pos COVID19 test result
a0_26|NA|presumed pos COVID19 result
a0_26|NA|presumed pos COVID test result
a0_26|NA|presumed pos COVID result
a0_26|NA|presumed pos for 2019 novel coronavirus
a0_26|NA|presumed pos for novel coronavirus
a0_26|NA|presumed pos for COVID 19
a0_26|NA|presumed pos for COVID19
a0_26|NA|presumed pos for COVID
a0_26|NA|presumed pos for 2019 novel coronavirus RNA
a0_26|NA|presumed pos for novel coronavirus RNA
a0_26|NA|presumed pos for COVID 19 RNA
a0_26|NA|presumed pos for COVID19 RNA
a0_27|NA|high temperatures
a0_27|NA|high temperature
a0_27|NA|fevered
a0_27|NA|fevering
a0_27|NA|feverish
a0_27|NA|fevers
a0_27|NA|fever
a0_27|NA|fièvre
a0_27|NA|fiver
a0_27|NA|feverin
a0_28|NA|CRISPR SARS-CoV-2 diagnostic test
a0_28|NA|CRISPR SARS-CoV-2 diagnostic testing
a0_28|NA|CRISPR SARS-CoV-2 diagnostic tests
a0_28|NA|CRISPR SARS-CoV-2 test
a0_28|NA|CRISPR SARS-CoV-2 testing
a0_28|NA|CRISPR SARS-CoV-2 tests
a0_28|NA|CRISPR SARS-CoV-2
a0_29|NA|COVID-19 spread
a0_29|NA|COVID-19 spreads
a0_29|NA|COVID-19 spreading
a0_29|NA|spread of COVID-19
a0_29|NA|COVID19 spread
a0_29|NA|COVID19 spreads
a0_29|NA|COVID19 spreading
a0_29|NA|spread of COVID19
a0_29|NA|COVID spread
a0_29|NA|COVID spreads
a0_29|NA|COVID spreading
a0_29|NA|spread of COVID
a0_29|NA|coronavirus spread
a0_29|NA|coronavirus spreads
a0_29|NA|coronavirus spreading
a0_29|NA|spread of coronavirus
a0_30|NA|COVID-toe
a0_30|NA|COVID-toes
a0_30|NA|sign of COVID-19
a0_30|NA|sign of COVID19
a0_30|NA|sign of COVID
a0_30|NA|chilblain-like lesions
a0_30|NA|chilblain-like lesion
a0_30|NA|chilblain-like
a0_30|NA|chilblain-like toe lesions
a0_30|NA|chilblain-like toe lesion
a0_31|NA|COVID-19 pandemic
a0_31|NA|COVID19 pandemic
a0_31|NA|COVID pandemic
a0_31|NA|coronavirus pandemic
a0_31|NA|COVID-19 outbreak
a0_31|NA|COVID19 outbreak
a0_31|NA|COVID outbreak
a0_31|NA|coronavirus outbreak
a0_31|NA|COVID-19 outbreaks
a0_31|NA|COVID19 outbreaks
a0_31|NA|COVID outbreaks
a0_31|NA|coronavirus outbreaks
a0_31|NA|outbreak of COVID-19
a0_31|NA|outbreak of COVID19
a0_31|NA|outbreak of COVID
a0_31|NA|outbreak of coronavirus
a0_31|NA|outbreaks of COVID-19
a0_31|NA|outbreaks of COVID19
a0_31|NA|outbreaks of COVID
a0_31|NA|outbreaks of coronavirus
a0_32|NA|COVID-19 pandemic
a0_32|NA|COVID19 pandemic
a0_32|NA|COVID pandemic
a0_32|NA|coronavirus pandemic
a0_32|NA|pandemic
a0_33|NA|non essential travel
a0_33|NA|non essential traveling
a0_33|NA|nonessential travel
a0_33|NA|nonessential traveling
a0_33|NA|traveling for non essential
a0_33|NA|traveling for nonessential
a0_33|NA|travel for non essential
a0_33|NA|travel for nonessential
a0_33|NA|travels for non essential
a0_33|NA|travels for nonessential
a0_33|NA|traveled for non essential
a0_33|NA|traveled for nonessential
a0_34|NA|COVID-19 signs and symptoms
a0_34|NA|signs and symptoms of COVID-19
a0_34|NA|COVID19 signs and symptoms
a0_34|NA|signs and symptoms of COVID19
a0_34|NA|COVID signs and symptoms
a0_34|NA|signs and symptoms of COVID
a0_34|NA|coronavirus signs and symptoms
a0_34|NA|signs and symptoms of coronavirus
a0_34|NA|signs and symptoms of the coronavirus
a0_34|NA|novel signs and symptoms
a0_34|NA|signs and symptoms of novel
a0_34|NA|signs and symptoms of the novel
a0_35|NA|dialyzability
a0_35|NA|dialyzabilities
a0_35|NA|dialysability
a0_35|NA|dialysabilities
a0_35|NA|dialysers
a0_35|NA|dialyser
a0_35|NA|dialysis solution
a0_35|NA|dialytic
a0_35|NA|dialyzers
a0_35|NA|dialyzer
a0_35|NA|dialysate
a0_35|NA|dialysis
a0_35|NA|dialyzable
a0_35|NA|dialyzing
a0_35|NA|dialyzes
a0_35|NA|dialyzed
a0_35|NA|dialyze
a0_35|NA|dialisys
a0_35|NA|dialyses
a0_35|NA|diaylisis
a0_35|NA|dialysi
a0_35|NA|dyalysis
a0_35|NA|dialisis
a0_35|NA|dialyisis
a0_35|NA|dialys
a0_35|NA|dialysus
a0_35|NA|diayliss
a0_35|NA|diaslysis
a0_35|NA|dailysis
a0_35|NA|diakysis
a0_35|NA|dialuysis
a0_35|NA|dialze
a0_35|NA|sialysis
a0_35|NA|dialysiys
a0_35|NA|dizlysis
a0_35|NA|ialysis
a0_35|NA|dialyz
a0_35|NA|dialyziable
a0_35|NA|dialytsis
a0_35|NA|dialystate
a0_35|NA|dialyzied
a0_35|NA|didalysis
a0_35|NA|diolysis
a0_35|NA|dialyzng
a0_35|NA|dialisate
a0_35|NA|dialyzier
a0_35|NA|ialyze
a0_35|NA|dialysiate
a0_35|NA|dialyzyed
a0_35|NA|dialysat
a0_35|NA|dialyyzing
a0_35|NA|cialyzer
a0_35|NA|dialyzsis
a0_35|NA|dialying
a0_35|NA|dlalysis
a0_35|NA|diablysis
a0_35|NA|dizlyzes
a0_35|NA|dializing
a0_35|NA|sialyzing
a0_35|NA|dialasis
a0_35|NA|sialyzed
a0_35|NA|dalysis
a0_35|NA|dialytics
a0_35|NA|doialysis
a0_35|NA|dialyizes
a0_35|NA|diualyzing
a0_35|NA|dialzying
a0_35|NA|dialyized
a0_35|NA|cialysis
a0_35|NA|dailyzing
a0_35|NA|dailyze
a0_35|NA|dialyssis
a0_35|NA|dialyste
a0_35|NA|dialysies
a0_35|NA|diealysis
a0_35|NA|dialyssi
a0_35|NA|dialyitic
a0_35|NA|dailysate
a0_35|NA|hdialysis
a0_35|NA|dialaysate
a0_35|NA|diazlyzed
a0_35|NA|dialkysis
a0_35|NA|ialyzing
a0_35|NA|dialyyzed
a0_35|NA|dialbysis
a0_35|NA|dialzing
a0_35|NA|dialyxing
a0_35|NA|dialysatem
a0_35|NA|dialylsate
a0_35|NA|dialysatel
a0_35|NA|adialysis
a0_35|NA|dialysates
a0_35|NA|dialasate
a0_35|NA|dialyvate
a0_35|NA|dialysaste
a0_35|NA|dialyusate
a0_35|NA|dilysate
a0_35|NA|qdialysate
a0_35|NA|dualysis
a0_35|NA|diayzer
a0_35|NA|duialysis
a0_35|NA|doialyze
a0_35|NA|dislyze
a0_35|NA|ialysate
a0_35|NA|dislysis
a0_35|NA|dialysated
a0_35|NA|dialyusis
a0_35|NA|dialoysis
a0_35|NA|dialyezd
a0_35|NA|dialystae
a0_35|NA|dializers
a0_35|NA|dialysed
a0_35|NA|dialsate
a0_35|NA|tdialysis
a0_35|NA|fdialysis
a0_35|NA|deialysis
a0_35|NA|dianlysis
a0_35|NA|dialyysis
a0_35|NA|disalysate
a0_35|NA|dialsyate
a0_35|NA|dialyaste
a0_35|NA|ndialysis
a0_35|NA|dialayzed
a0_35|NA|dialyzate
a0_35|NA|dialytis
a0_35|NA|diallysate
a0_35|NA|dioalysis
a0_35|NA|dialysyis
a0_35|NA|dialye
a0_35|NA|dislyzes
a0_35|NA|diayzing
a0_35|NA|dialyzzed
a0_35|NA|diaysis
a0_35|NA|qdialysis
a0_35|NA|diahysis
a0_35|NA|dialylzing
a0_35|NA|dialyuzed
a0_35|NA|diaysate
a0_35|NA|dialysiis
a0_35|NA|dialyiss
a0_35|NA|dislysate
a0_35|NA|dialylze
a0_35|NA|dialyate
a0_35|NA|dialysis1
a0_35|NA|dialylsis
a0_35|NA|dializes
a0_35|NA|dializer
a0_35|NA|dialysis2
a0_35|NA|tialysis
a0_35|NA|rialysis
a0_35|NA|dialyaed
a0_35|NA|dilayzed
a0_35|NA|dialzyzed
a0_35|NA|dialyslate
a0_35|NA|gdialysis
a0_35|NA|dilayzing
a0_35|NA|dialyizing
a0_35|NA|diallysis
a0_35|NA|dilalyze
a0_35|NA|dialized
a0_35|NA|dialyasis
a0_35|NA|dialyizable
a0_35|NA|dilaytic
a0_35|NA|dialyisate
a0_35|NA|dialzyzes
a0_35|NA|dialaysis
a0_35|NA|dialyzeer
a0_35|NA|dialysze
a0_35|NA|dilaysate
a0_35|NA|diaylysis
a0_35|NA|dialhysis
a0_35|NA|doalyzing
a0_35|NA|dialyzine
a0_35|NA|dialysys
a0_35|NA|dialysic
a0_35|NA|dialysid
a0_35|NA|dialysie
a0_35|NA|dialzye
a0_35|NA|dialysia
a0_35|NA|dialysil
a0_35|NA|dializable
a0_35|NA|dialysios
a0_35|NA|dilaysis
a0_35|NA|dialize
a0_35|NA|diaclysis
a0_35|NA|dialyzying
a0_35|NA|dialsysate
a0_35|NA|dialyazes
a0_35|NA|disalysis
a0_35|NA|dialylzed
a0_35|NA|diaylze
a0_35|NA|dilayze
a0_35|NA|dialyazed
a0_35|NA|dalysate
a0_35|NA|dialylate
a0_35|NA|dialyis
a0_35|NA|ddialysis
a0_35|NA|diayzed
a0_35|NA|dialysins
a0_35|NA|diaytic
a0_35|NA|diaiysis
a0_35|NA|dalyze
a0_35|NA|dailytic
a0_35|NA|dialyzi
a0_35|NA|dilalysis
a0_35|NA|dialyzin
a0_35|NA|dixlyze
a0_35|NA|odialysis
a0_35|NA|dialysing
a0_35|NA|diaylyzes
a0_35|NA|dailyzer
a0_35|NA|dailyzed
a0_35|NA|dialsysis
a0_35|NA|dialosis
a0_35|NA|dialyzis
a0_35|NA|diaylzed
a0_35|NA|dialyzzd
a0_35|NA|diapysis
a0_35|NA|dilayzes
a0_35|NA|dialyzie
a0_35|NA|dialaze
a0_35|NA|dialyxed
a0_35|NA|dialyzig
a0_35|NA|dxalyze
a0_35|NA|diaylzes
a0_35|NA|dialyziing
a0_35|NA|dialysius
a0_35|NA|dialusate
a0_35|NA|dialysls
a0_35|NA|dialyhsis
a0_35|NA|dialzyes
a0_35|NA|diaoysis
a0_35|NA|dialyasate
a0_35|NA|dialyss
a0_35|NA|dialzed
a0_35|NA|dilysis
a0_35|NA|dialyszing
a0_35|NA|dialsyze
a0_35|NA|dialsyis
a0_35|NA|dialzer
a0_35|NA|doialyzed
a0_35|NA|dialynate
a0_35|NA|mdialysis
a0_35|NA|dialyable
a0_35|NA|diialyzed
a0_35|NA|dilalyzed
a0_35|NA|dialzyed
a0_35|NA|dialyti
a0_35|NA|dialysyte
a0_35|NA|dialzes
a0_35|NA|dialyte
a0_35|NA|dialyszer
a0_35|NA|diaplysis
a0_35|NA|pdialysis
a0_35|NA|dialyctic
a0_35|NA|dialiysis
a0_35|NA|dsialysis
a0_35|NA|dialystis
a0_35|NA|dialusis
a0_35|NA|ialyzable
a0_35|NA|dialysite
a0_35|NA|dialyyze
a0_35|NA|idalysis
a0_35|NA|dialyslis
a0_35|NA|dialyszed
a0_35|NA|dialyais
a0_35|NA|dialyaze
a0_35|NA|dialysdis
a0_35|NA|dialystic
a0_35|NA|diaylsate
a0_35|NA|dialysisz
a0_35|NA|dialysist
a0_35|NA|dialyize
a0_35|NA|dilyzed
a0_35|NA|dialysiss
a0_35|NA|doalysis
a0_35|NA|dialysisr
a0_35|NA|dialysism
a0_35|NA|dialysisl
a0_35|NA|diialysis
a0_35|NA|dialysisn
a0_35|NA|dialsis
a0_35|NA|ialyzed
a0_35|NA|dialysise
a0_35|NA|diasysis
a0_35|NA|dialyed
a0_35|NA|daalysis
a0_35|NA|dialysisf
a0_35|NA|diaylzing
a0_35|NA|dialysisa
a0_35|NA|dilyzes
a0_35|NA|dialyes
a0_35|NA|dialysable
a0_35|NA|ialytic
a0_35|NA|daialysis
a0_35|NA|dilyze
a0_35|NA|eialysis
a0_35|NA|dialysuis
a0_35|NA|dialysias
a0_35|NA|rdialyzed
a0_35|NA|dialyssate
a0_35|NA|diayze
a0_35|NA|mialysis
a0_35|NA|dialyzede
a0_35|NA|dialysis8
a0_35|NA|dialysos
a0_35|NA|ialyzes
a0_35|NA|ialyzer
a0_35|NA|dialysis4
a0_35|NA|dialysis6
a0_35|NA|diualysis
a0_35|NA|dyalisate
a0_35|NA|dyalizer
a0_35|NA|dyalizers
a0_35|NA|diaalysis
a0_36|NA|fever rose
a0_36|NA|temperature was raised
a0_36|NA|temperature is raised
a0_36|NA|temperature raised
a0_36|NA|temperatures are raised
a0_36|NA|temperature were raised
a0_36|NA|raised temperature
a0_36|NA|raised temperatures
a0_36|NA|body temperature was raised
a0_36|NA|body temperature is raised
a0_36|NA|body temperature raised
a0_36|NA|body temperatures are raised
a0_36|NA|body temperature were raised
a0_36|NA|raised body temperature
a0_36|NA|raised body temperatures
a0_36|NA|temp was raised
a0_36|NA|temp is raised
a0_36|NA|temp raised
a0_36|NA|temps are raised
a0_36|NA|temp were raised
a0_36|NA|raised temp
a0_36|NA|raised temps
a0_36|NA|body temp was raised
a0_36|NA|body temp is raised
a0_36|NA|body temp raised
a0_36|NA|body temps are raised
a0_36|NA|body temp were raised
a0_36|NA|raised body temp
a0_36|NA|raised body temps
a0_36|NA|increase in body temperature
a0_36|NA|spiking a fever
a0_36|NA|spiked a fever
a0_36|NA|spikes a fever
a0_36|NA|spike a fever
a0_36|NA|fever spikes
a0_36|NA|fever spike
a0_36|NA|spiking fevers
a0_36|NA|spiking fever
a0_36|NA|spiked fevers
a0_36|NA|spiked fever
a0_36|NA|spikes fevers
a0_36|NA|spikes fever
a0_36|NA|spike fevers
a0_36|NA|spike fever
a0_36|NA|febrility
a0_36|NA|febrile
a0_36|NA|feverishness
a0_36|NA|feverish
a0_36|NA|fevers
a0_36|NA|fever
a0_36|NA|temperatures
a0_36|NA|temperature
a0_36|NA|temps
a0_36|NA|temp
a0_36|NA|pyretics
a0_36|NA|pyretic
a0_36|NA|pyrexial
a0_36|NA|pyrexic
a0_36|NA|hyper-pyrexial
a0_36|NA|hyper-pyrexia
a0_36|NA|hyper-pyrexic
a0_36|NA|hyperpyrexial
a0_36|NA|hyperpyrexia
a0_36|NA|hyperpyrexic
a0_36|NA|pyrexia
a0_36|NA|T-max
a0_36|NA|Tmax
a0_36|NA|Tm
a0_36|NA|burning up
a0_36|NA|feeling hot
a0_36|NA|feels hot
a0_36|NA|felt hot
a0_36|NA|feel hot
a0_36|NA|forehead feels hot
a0_36|NA|forehead felt hot
a0_36|NA|forehead was feeling hot
a0_36|NA|hot to the touch
a0_36|NA|hot to touch
a0_36|NA|feeling warm
a0_36|NA|feels warm
a0_36|NA|felt warm
a0_36|NA|feel warm
a0_36|NA|forehead feels warm
a0_36|NA|forehead felt warm
a0_36|NA|forehead was feeling warm
a0_36|NA|warm to the touch
a0_36|NA|warm to touch
a0_36|NA|febirle
a0_36|NA|fevr
a0_36|NA|fevor
a0_36|NA|feberile
a0_36|NA|feveer
a0_36|NA|feverk
a0_37|NA|school closures
a0_37|NA|school closure
a0_37|NA|schools are closed
a0_37|NA|schools closed
a0_37|NA|school is closed
a0_37|NA|school closed
a0_37|NA|schools are closing
a0_37|NA|schools closing
a0_37|NA|school is closing
a0_37|NA|school closing
a0_37|NA|school closings
a0_37|NA|closing the schools
a0_37|NA|closing the school
a0_37|NA|closing schools
a0_37|NA|closing school
a0_37|NA|closed the schools
a0_37|NA|closed the school
a0_37|NA|closed schools
a0_37|NA|closed school
a0_37|NA|closes the schools
a0_37|NA|closes the school
a0_37|NA|closes schools
a0_37|NA|closes school
a0_37|NA|close the schools
a0_37|NA|close the school
a0_37|NA|close schools
a0_37|NA|close school
a0_38|NA|COVID-19 tent
a0_38|NA|COVID-19 tents
a0_38|NA|COVID19 tent
a0_38|NA|COVID19 tents
a0_38|NA|COVID tent
a0_38|NA|COVID tents
a0_38|NA|coronavirus tent
a0_38|NA|coronavirus tents
a0_39|NA|COVID-19 infection
a0_39|NA|COVID-19
a0_39|NA|2019-nCoV acute respiratory disease
a0_39|NA|U07.1
a0_40|NA|first human trial
a0_40|NA|first human trials
a0_40|NA|human trial
a0_40|NA|human trials
a0_40|NA|first trial in humans
a0_40|NA|first trials in humans
a0_40|NA|trial in humans
a0_40|NA|trials in humans
a0_41|NA|toxicity of hydroxychloroquine
a0_41|NA|toxicities of hydroxychloroquine
a0_41|NA|hydroxychloroquine toxicity
a0_41|NA|hydroxychloroquine toxicities
a0_41|NA|hydroxychloroquine tox
a0_41|NA|toxicity of HCQ
a0_41|NA|toxicities of HCQ
a0_41|NA|HCQ toxicity
a0_41|NA|HCQ toxicities
a0_41|NA|HCQ tox
a0_41|NA|toxicity of Plaquenil
a0_41|NA|toxicities of Plaquenil
a0_41|NA|Plaquenil toxicity
a0_41|NA|Plaquenil toxicities
a0_41|NA|Plaquenil tox
a0_41|NA|intoxicated by HCQ
a0_41|NA|intoxicated from HCQ
a0_41|NA|intoxication from HCQ
a0_41|NA|intoxications from HCQ
a0_41|NA|poisoned by HCQ
a0_41|NA|poisoning from HCQ
a0_41|NA|HCQ-induced intoxication
a0_41|NA|HCQ-induced poisoning
a0_41|NA|HCQ-induced toxicities
a0_41|NA|HCQ intoxications
a0_41|NA|HCQ intoxication
a0_41|NA|HCQ poisonings
a0_41|NA|intoxicated by hydroxychloroquine
a0_41|NA|intoxicated from hydroxychloroquine
a0_41|NA|intoxication from hydroxychloroquine
a0_41|NA|intoxications from hydroxychloroquine
a0_41|NA|poisoned by hydroxychloroquine
a0_41|NA|poisoning from hydroxychloroquine
a0_41|NA|hydroxychloroquine-induced intoxication
a0_41|NA|hydroxychloroquine-induced poisoning
a0_41|NA|hydroxychloroquine-induced toxicities
a0_41|NA|hydroxychloroquine intoxications
a0_41|NA|hydroxychloroquine intoxication
a0_41|NA|hydroxychloroquine poisonings
a0_41|NA|toxic side effects of hydroxychloroquine
a0_41|NA|toxic side effect of hydroxychloroquine
a0_41|NA|toxic effects of hydroxychloroquine
a0_41|NA|toxic effect of hydroxychloroquine
a0_41|NA|side effects of hydroxychloroquine
a0_41|NA|side effect of hydroxychloroquine
a0_41|NA|hydroxychloroquine side effects
a0_41|NA|hydroxychloroquine side effect
a0_41|NA|hydroxychloroquine poisoning
a0_41|NA|hydroxychloroquine-induced toxicity
a0_41|NA|toxic side effects of HCQ
a0_41|NA|toxic side effect of HCQ
a0_41|NA|toxic effects of HCQ
a0_41|NA|toxic effect of HCQ
a0_41|NA|side effects of HCQ
a0_41|NA|side effect of HCQ
a0_41|NA|HCQ side effects
a0_41|NA|HCQ side effect
a0_41|NA|HCQ poisoning
a0_41|NA|HCQ-induced toxicity
a0_41|NA|intoxicated by Plaquenil
a0_41|NA|intoxicated from Plaquenil
a0_41|NA|intoxication from Plaquenil
a0_41|NA|intoxications from Plaquenil
a0_41|NA|poisoned by Plaquenil
a0_41|NA|poisoning from Plaquenil
a0_41|NA|Plaquenil-induced intoxication
a0_41|NA|Plaquenil-induced poisoning
a0_41|NA|Plaquenil-induced toxicities
a0_41|NA|Plaquenil intoxications
a0_41|NA|Plaquenil intoxication
a0_41|NA|Plaquenil poisonings
a0_41|NA|toxic side effects of Plaquenil
a0_41|NA|toxic side effect of Plaquenil
a0_41|NA|toxic effects of Plaquenil
a0_41|NA|toxic effect of Plaquenil
a0_41|NA|side effects of Plaquenil
a0_41|NA|side effect of Plaquenil
a0_41|NA|Plaquenil side effects
a0_41|NA|Plaquenil side effect
a0_41|NA|Plaquenil poisoning
a0_41|NA|Plaquenil-induced toxicity
a0_41|NA|Plaquenil
a0_41|NA|HCQ
a0_41|NA|hydroxychloroquine
a0_42|NA|COVID-19 cases
a0_42|NA|COVID-19 case
a0_42|NA|COVID19 cases
a0_42|NA|COVID19 case
a0_42|NA|COVID cases
a0_42|NA|COVID case
a0_42|NA|coronavirus cases
a0_42|NA|coronavirus case
a0_42|NA|cases of COVID-19
a0_42|NA|cases of COVID19
a0_42|NA|cases of COVID
a0_42|NA|cases of coronavirus
a0_42|NA|case of COVID-19
a0_42|NA|case of COVID19
a0_42|NA|case of COVID
a0_42|NA|case of coronavirus
a0_42|NA|diagnosed with COVID-19
a0_42|NA|diagnosed with COVID19
a0_42|NA|diagnosed with COVID
a0_42|NA|diagnosed with coronavirus
a0_42|NA|COVID-19 diagnosis
a0_42|NA|COVID-19 diagnoses
a0_42|NA|COVID19 diagnosis
a0_42|NA|COVID19 diagnoses
a0_42|NA|COVID diagnosis
a0_42|NA|COVID diagnoses
a0_42|NA|coronavirus diagnosis
a0_42|NA|coronavirus diagnoses
a0_42|NA|diagnosis of COVID-19
a0_42|NA|diagnosis of COVID19
a0_42|NA|diagnosis of COVID
a0_42|NA|COVID-19 patients
a0_42|NA|COVID-19 patient
a0_42|NA|COVID19 patients
a0_42|NA|COVID19 patient
a0_42|NA|COVID patient
a0_42|NA|COVID patients
a0_42|NA|coronavirus patients
a0_42|NA|coronavirus patient
a0_42|NA|patients with COVID-19
a0_42|NA|patients with COVID19
a0_42|NA|patients with COVID
a0_42|NA|patients with coronavirus
a0_42|NA|patients diagnosed with COVID-19
a0_42|NA|patients diagnosed with COVID19
a0_42|NA|patients diagnosed with COVID
a0_42|NA|patients diagnosed with coronavirus
a0_42|NA|patients with a diagnosis of COVID-19
a0_42|NA|patients with diagnosis of COVID-19
a0_42|NA|patients with a diagnosis of COVID19
a0_42|NA|patients with diagnosis of COVID19
a0_42|NA|patients with a diagnosis of COVID
a0_42|NA|patients with diagnosis of COVID
a0_42|NA|patients with a diagnosis of coronavirus
a0_42|NA|patients with diagnosis of coronavirus
a0_42|NA|patient with COVID-19
a0_42|NA|patient with COVID19
a0_42|NA|patient with COVID
a0_42|NA|patient with coronavirus
a0_42|NA|patient diagnosed with COVID-19
a0_42|NA|patient diagnosed with COVID19
a0_42|NA|patient diagnosed with COVID
a0_42|NA|patient diagnosed with coronavirus
a0_42|NA|patient with a diagnosis of COVID-19
a0_42|NA|patient with diagnosis of COVID-19
a0_42|NA|patient with a diagnosis of COVID19
a0_42|NA|patient with diagnosis of COVID19
a0_42|NA|patient with a diagnosis of COVID
a0_42|NA|patient with diagnosis of COVID
a0_42|NA|patient with a diagnosis of coronavirus
a0_42|NA|patient with diagnosis of coronavirus
a0_43|NA|COVID-19 pandemic
a0_43|NA|COVID19 pandemic
a0_43|NA|COVID pandemic
a0_43|NA|coronavirus pandemic
a0_45|NA|pneumonia due to 2019 novel coronavirus
a0_45|NA|pneumonia due to 2019 coronavirus
a0_45|NA|pneumonia due to coronavirus
a0_45|NA|pneumonia due to COVID-19
a0_45|NA|pneumonia due to COVID19
a0_45|NA|pneumonia due to COVID
a0_45|NA|pneumonia secondary to 2019 novel coronavirus
a0_45|NA|pneumonia secondary to 2019 coronavirus
a0_45|NA|pneumonia secondary to coronavirus
a0_45|NA|pneumonia secondary to COVID-19
a0_45|NA|pneumonia secondary to COVID19
a0_45|NA|pneumonia secondary to COVID
a0_45|NA|2019 novel coronavirus pneumonia
a0_45|NA|novel coronavirus pneumonia
a0_45|NA|2019 coronavirus pneumonia
a0_45|NA|coronavirus pneumonia
a0_45|NA|COVID-19 pneumonia
a0_45|NA|COVID19 pneumonia
a0_45|NA|COVID pneumonia
a0_45|NA|2019 novel coronavirus with pneumonia
a0_45|NA|2019 coronavirus with pneumonia
a0_45|NA|coronavirus with pneumonia
a0_45|NA|COVID-19 with pneumonia
a0_45|NA|COVID19 with pneumonia
a0_45|NA|COVID with pneumonia
a0_45|NA|2019 novel coronavirus complicated by pneumonia
a0_45|NA|2019 coronavirus complicated by pneumonia
a0_45|NA|coronavirus complicated by pneumonia
a0_45|NA|COVID-19 complicated by pneumonia
a0_45|NA|COVID19 complicated by pneumonia
a0_45|NA|COVID complicated by pneumonia
a0_45|NA|PNA due to 2019 novel coronavirus
a0_45|NA|PNA due to 2019 coronavirus
a0_45|NA|PNA due to coronavirus
a0_45|NA|PNA due to COVID-19
a0_45|NA|PNA due to COVID19
a0_45|NA|PNA due to COVID
a0_45|NA|PNA secondary to 2019 novel coronavirus
a0_45|NA|PNA secondary to 2019 coronavirus
a0_45|NA|PNA secondary to coronavirus
a0_45|NA|PNA secondary to COVID-19
a0_45|NA|PNA secondary to COVID19
a0_45|NA|PNA secondary to COVID
a0_45|NA|2019 novel coronavirus PNA
a0_45|NA|2019 coronavirus PNA
a0_45|NA|coronavirus PNA
a0_45|NA|COVID-19 PNA
a0_45|NA|COVID19 PNA
a0_45|NA|COVID PNA
a0_45|NA|2019 novel coronavirus with PNA
a0_45|NA|2019 coronavirus with PNA
a0_45|NA|coronavirus with PNA
a0_45|NA|COVID-19 with PNA
a0_45|NA|COVID19 with PNA
a0_45|NA|COVID with PNA
a0_45|NA|2019 novel coronavirus complicated by PNA
a0_45|NA|2019 coronavirus complicated by PNA
a0_45|NA|coronavirus complicated by PNA
a0_45|NA|COVID-19 complicated by PNA
a0_45|NA|COVID19 complicated by PNA
a0_45|NA|COVID complicated by PNA
a0_46|NA|first human drug trial
a0_46|NA|first human drug trials
a0_46|NA|first human trial
a0_46|NA|first human trials
a0_46|NA|first drug trial in humans
a0_46|NA|first drug trials in humans
a0_47|NA|COVID-19 test kits
a0_47|NA|COVID-19 test kit
a0_47|NA|test kit for COVID-19
a0_47|NA|test kits for COVID-19
a0_47|NA|COVID-19 testing kits
a0_47|NA|COVID-19 testing kit
a0_47|NA|testing kit for COVID-19
a0_47|NA|testing kits for COVID-19
a0_47|NA|COVID19 test kits
a0_47|NA|COVID19 test kit
a0_47|NA|test kit for COVID19
a0_47|NA|test kits for COVID19
a0_47|NA|COVID19 testing kits
a0_47|NA|COVID19 testing kit
a0_47|NA|testing kit for COVID19
a0_47|NA|testing kits for COVID19
a0_47|NA|coronavirus test kits
a0_47|NA|coronavirus test kit
a0_47|NA|test kit for coronavirus
a0_47|NA|test kits for coronavirus
a0_47|NA|coronavirus testing kits
a0_47|NA|coronavirus testing kit
a0_47|NA|testing kit for coronavirus
a0_47|NA|testing kits for coronavirus
a0_47|NA|COVID test kits
a0_47|NA|COVID test kit
a0_47|NA|test kit for COVID
a0_47|NA|test kits for COVID
a0_47|NA|COVID testing kits
a0_47|NA|COVID testing kit
a0_47|NA|testing kit for COVID
a0_47|NA|testing kits for COVID
a0_48|NA|practicing social distancing
a0_48|NA|practiced social distancing
a0_48|NA|practices social distancing
a0_48|NA|practice social distancing
a0_48|NA|social distancing
a0_49|NA|first human vaccine trial
a0_49|NA|first human vaccine trials
a0_49|NA|first human trial
a0_49|NA|first human trials
a0_49|NA|first vaccine trial in humans
a0_49|NA|first vaccine trials in humans
a0_50|NA|non-COVID-19
a0_50|NA|non-COVID19
a0_50|NA|non-COVID
a0_50|NA|non-coronavirus
a0_50|NA|nonCOVID-19
a0_50|NA|nonCOVID19
a0_50|NA|nonCOVID
a0_50|NA|noncoronavirus
a0_50|NA|not COVID-19
a0_50|NA|not COVID19
a0_50|NA|not COVID
a0_50|NA|not coronavirus
a0_50|NA|not the coronavirus
a0_50|NA|not the novel coronavirus
a0_51|NA|hydroxychloroquine
a0_51|NA|Hidroxicloroquina
a0_51|NA|Hydroxychlorochin
a0_51|NA|Hydroxychloroguine
a0_51|NA|Hydroxychloroquinum
a0_51|NA|Idrossiclorochina
a0_51|NA|Oxichlorochine
a0_51|NA|Oxichlorochinum
a0_51|NA|Oxichloroquine
a0_51|NA|Oxychlorochin
a0_51|NA|Oxychloroquine
a0_51|NA|Polirreumin
a0_51|NA|Quensyl
a0_51|NA|WIN 1258
a0_51|NA|WIN1258
a0_52|NA|confirmed positive coronavirus
a0_52|NA|confirmed positive for coronavirus
a0_52|NA|confirmed pos coronavirus
a0_52|NA|confirmed pos for coronavirus
a0_52|NA|confirmed coronavirus
a0_52|NA|coronavirus testing was positive
a0_52|NA|coronavirus test was positive
a0_52|NA|coronavirus testing was pos
a0_52|NA|coronavirus test was pos
a0_52|NA|coronavirus testing is positive
a0_52|NA|coronavirus test is positive
a0_52|NA|coronavirus testing is pos
a0_52|NA|coronavirus test is pos
a0_52|NA|tested positive coronavirus
a0_52|NA|tested positive for coronavirus
a0_52|NA|tested pos coronavirus
a0_52|NA|tested pos for coronavirus
a0_52|NA|tested positive for the coronavirus
a0_52|NA|tested positive for the novel coronavirus
a0_52|NA|tested pos for the coronavirus
a0_52|NA|tested pos for the novel coronavirus
a0_52|NA|confirmed positive COVID19
a0_52|NA|confirmed positive COVID-19
a0_52|NA|confirmed positive for COVID19
a0_52|NA|confirmed positive for COVID-19
a0_52|NA|confirmed pos COVID19
a0_52|NA|confirmed pos COVID-19
a0_52|NA|confirmed pos for COVID19
a0_52|NA|confirmed pos for COVID-19
a0_52|NA|confirmed COVID19
a0_52|NA|confirmed COVID-19
a0_52|NA|COVID19 testing was positive
a0_52|NA|COVID19 test was positive
a0_52|NA|COVID-19 testing was positive
a0_52|NA|COVID-19 test was positive
a0_52|NA|COVID19 testing was pos
a0_52|NA|COVID19 test was pos
a0_52|NA|COVID-19 testing was pos
a0_52|NA|COVID-19 test was pos
a0_52|NA|COVID19 testing is positive
a0_52|NA|COVID19 test is positive
a0_52|NA|COVID-19 testing is positive
a0_52|NA|COVID-19 test is positive
a0_52|NA|COVID19 testing is pos
a0_52|NA|COVID19 test is pos
a0_52|NA|COVID-19 testing is pos
a0_52|NA|COVID-19 test is pos
a0_52|NA|tested positive COVID19
a0_52|NA|tested positive COVID-19
a0_52|NA|tested positive for COVID19
a0_52|NA|tested positive for COVID-19
a0_52|NA|tested pos COVID19
a0_52|NA|tested pos COVID-19
a0_52|NA|tested pos for COVID19
a0_52|NA|tested pos for COVID-19
a0_52|NA|COVID19 test positive
a0_52|NA|COVID 19 test positive
a0_52|NA|coronavirus test positive
a0_52|NA|COVID19 test pos
a0_52|NA|COVID 19 test pos
a0_52|NA|coronavirus test pos
a0_52|NA|COVID 19 positive
a0_52|NA|COVID19 positive
a0_52|NA|COVID positive
a0_52|NA|2019 novel coronavirus positive
a0_52|NA|COVID 19 PCR positive for 2019 novel coronavirus
a0_52|NA|PCR positive for 2019 novel coronavirus
a0_52|NA|PCR positive for novel coronavirus
a0_52|NA|PCR positive for COVID 19
a0_52|NA|PCR positive for COVID19
a0_52|NA|PCR positive for COVID
a0_52|NA|positive COVID 19 test result
a0_52|NA|positive COVID 19 result
a0_52|NA|positive COVID19 test result
a0_52|NA|positive COVID19 result
a0_52|NA|positive COVID test result
a0_52|NA|positive COVID result
a0_52|NA|positive for 2019 novel coronavirus
a0_52|NA|positive for novel coronavirus
a0_52|NA|positive for COVID 19
a0_52|NA|positive for COVID19
a0_52|NA|positive for COVID
a0_52|NA|positive for 2019 novel coronavirus RNA
a0_52|NA|positive for novel coronavirus RNA
a0_52|NA|positive for COVID 19 RNA
a0_52|NA|positive for COVID19 RNA
a0_52|NA|positive for COVID RNA
a0_52|NA|real time PCR positive for 2019 novel coronavirus
a0_52|NA|real time PCR positive for novel coronavirus
a0_52|NA|real time PCR positive for coronavirus
a0_52|NA|real time PCR positive for COVID 19
a0_52|NA|real time PCR positive for COVID19
a0_52|NA|real time PCR positive for COVID
a0_52|NA|COVID 19 pos
a0_52|NA|COVID19 pos
a0_52|NA|COVID pos
a0_52|NA|2019 novel coronavirus pos
a0_52|NA|COVID 19 PCR pos for 2019 novel coronavirus
a0_52|NA|PCR pos for 2019 novel coronavirus
a0_52|NA|PCR pos for novel coronavirus
a0_52|NA|PCR pos for COVID 19
a0_52|NA|PCR pos for COVID19
a0_52|NA|PCR pos for COVID
a0_52|NA|pos COVID 19 test result
a0_52|NA|pos COVID 19 result
a0_52|NA|pos COVID19 test result
a0_52|NA|pos COVID19 result
a0_52|NA|pos COVID test result
a0_52|NA|pos COVID result
a0_52|NA|pos for 2019 novel coronavirus
a0_52|NA|pos for novel coronavirus
a0_52|NA|pos for COVID 19
a0_52|NA|pos for COVID19
a0_52|NA|pos for COVID
a0_52|NA|pos for 2019 novel coronavirus RNA
a0_52|NA|pos for novel coronavirus RNA
a0_52|NA|pos for COVID 19 RNA
a0_52|NA|pos for COVID19 RNA
a0_52|NA|pos for COVID RNA
a0_52|NA|real time PCR pos for 2019 novel coronavirus
a0_52|NA|real time PCR pos for novel coronavirus
a0_52|NA|real time PCR pos for coronavirus
a0_52|NA|real time PCR pos for COVID 19
a0_52|NA|real time PCR pos for COVID19
a0_52|NA|real time PCR pos for COVID
a0_53|NA|COVID-19 symptoms
a0_53|NA|COVID-19 symptom
a0_53|NA|symptoms of COVID-19
a0_53|NA|symptom of COVID-19
a0_53|NA|COVID19 symptoms
a0_53|NA|COVID19 symptom
a0_53|NA|symptoms of COVID19
a0_53|NA|symptom of COVID19
a0_53|NA|COVID symptoms
a0_53|NA|COVID symptom
a0_53|NA|symptoms of COVID
a0_53|NA|symptom of COVID
a0_53|NA|coronavirus symptoms
a0_53|NA|coronavirus symptom
a0_53|NA|symptoms of coronavirus
a0_53|NA|symptom of coronavirus
a0_53|NA|symptoms of the coronavirus
a0_53|NA|symptom of the coronavirus
a0_53|NA|novel symptoms
a0_53|NA|novel symptom
a0_53|NA|symptoms of novel
a0_53|NA|symptom of novel
a0_53|NA|symptoms of the novel
a0_53|NA|symptom of the novel
a0_54|NA|oropharyngeal swabs
a0_54|NA|oropharyngeal swab
a0_54|NA|oropharyngeal sample
a0_54|NA|oropharyngeal samples
a0_54|NA|oropharyngeal sampling
a0_54|NA|oro-pharyngeal swabs
a0_54|NA|oro-pharyngeal swab
a0_54|NA|oro-pharyngeal sample
a0_54|NA|oro-pharyngeal samples
a0_54|NA|oro-pharyngeal sampling
a0_54|NA|oropharynx swabs
a0_54|NA|oropharynx swab
a0_54|NA|oropharynx sample
a0_54|NA|oropharynx samples
a0_54|NA|oropharynx sampling
a0_54|NA|oro-pharynx swabs
a0_54|NA|oro-pharynx swab
a0_54|NA|oro-pharynx sample
a0_54|NA|oro-pharynx samples
a0_54|NA|oro-pharynx sampling
a0_54|NA|OP swabs
a0_54|NA|OP swab
a0_54|NA|OP sample
a0_54|NA|OP samples
a0_54|NA|OP sampling
a0_54|NA|swabbing the OP
a0_54|NA|swabbing the oro-pharynx
a0_54|NA|swabbing the oropharynx
a0_54|NA|swabbed the OP
a0_54|NA|swabbed the oro-pharynx
a0_54|NA|swabbed the oropharynx
a0_54|NA|swabs the OP
a0_54|NA|swabs the oro-pharynx
a0_54|NA|swabs the oropharynx
a0_54|NA|swab the OP
a0_54|NA|swab the oro-pharynx
a0_54|NA|swab the oropharynx
a0_54|NA|samples from the OP
a0_54|NA|sample from the OP
a0_54|NA|samples from OP
a0_54|NA|sample from OP
a0_54|NA|samples from the oropharynx
a0_54|NA|sample from the oropharynx
a0_54|NA|samples from oropharynx
a0_54|NA|sample from oropharynx
a0_54|NA|samples from the oro-pharynx
a0_54|NA|sample from the oro-pharynx
a0_54|NA|samples from oro-pharynx
a0_54|NA|sample from oro-pharynx
a0_54|NA|sampling the OP
a0_54|NA|sampled the OP
a0_54|NA|samples the OP
a0_54|NA|sample the OP
a0_54|NA|sampling the oropharynx
a0_54|NA|sampled the oropharynx
a0_54|NA|samples the oropharynx
a0_54|NA|sample the oropharynx
a0_54|NA|sampling the oro-pharynx
a0_54|NA|sampled the oro-pharynx
a0_54|NA|samples the oro-pharynx
a0_54|NA|sample the oro-pharynx
a0_55|NA|hydroxychloroquine
a0_55|NA|hydrossicloroquine
a0_55|NA|hydroxicloroquine
a0_55|NA|hydroxychlorochine
a0_55|NA|hydroxycloroquine
a0_55|NA|hydryxychloroquine
a0_55|NA|hydroxyxchloroquine
a0_55|NA|lhydroxychloroquine
a0_55|NA|hydroxychloroquinr
a0_55|NA|hydroxychloroquinne
a0_55|NA|hydropychloroquine
a0_55|NA|hydrdoxychloroquine
a0_55|NA|hydroxychloroqune
a0_55|NA|hydroxychloroquinw
a0_55|NA|hydroxychlorofuine
a0_55|NA|hydroxychloruquine
a0_55|NA|hydroxyxhloroquine
a0_55|NA|hydroxychloroquire
a0_55|NA|hydrozychloroquine
a0_55|NA|hydroyxychloroquine
a0_55|NA|hydroxychloroqiune
a0_55|NA|hydroychloroquine
a0_55|NA|hydroxycholoroquine
a0_55|NA|hydroxychloriquine
a0_55|NA|hydroxychloroquinet
a0_55|NA|hydroxychloroquinn
a0_55|NA|hydroxychloroqine
a0_55|NA|hydroxychlorozuine
a0_55|NA|hydrxychloroquine
a0_55|NA|hydroxichloroquine
a0_55|NA|hydroxychlorpquine
a0_55|NA|hydroxychloroquin
a0_55|NA|hydoxychloroquine
a0_55|NA|hydryoxychloroquine
a0_55|NA|hydroxychloroquien
a0_55|NA|hydroxychloroquie
a0_55|NA|hydroxhchloroquine
a0_55|NA|hydcroxychloroquine
a0_55|NA|hydroxychloraquine
a0_55|NA|dydroxychloroquine
a0_55|NA|hydtoxychloroquine
a0_55|NA|hydroxuchloroquine
a0_55|NA|hydroxyzhloroquine
a0_55|NA|hydroxychloroquiine
a0_55|NA|hydroxrychloroquine
a0_55|NA|hydroxchloroquine
a0_55|NA|hydroxychlorouqine
a0_55|NA|hydroxoychloroquine
a0_55|NA|hytroxychloroquine
a0_55|NA|hydroxychkoroquine
a0_55|NA|hydroyxchloroquine
a0_55|NA|hydroxycholroquine
a0_55|NA|hydroxyhloroquine
a0_55|NA|hydroxychloroquince
a0_55|NA|hyroxychloroquine
a0_55|NA|hdroxychloroquine
a0_55|NA|hydroxytchloroquine
a0_55|NA|ydroxychloroquine
a0_55|NA|hydroxylchloroquine
a0_55|NA|hyrdroxychloroquine
a0_55|NA|hydrocychloroquine
a0_55|NA|hydroxychlroquine
a0_55|NA|hydrooxychloroquine
a0_55|NA|hydroxcychloroquine
a0_55|NA|hdyroxychloroquine
a0_55|NA|hyrdoxychloroquine
a0_55|NA|hydroxzchloroquine
a0_55|NA|hhydroxychloroquine
a0_55|NA|hycroxychloroquine
a0_55|NA|hyxdroxychloroquine
a0_55|NA|hydroxychloloquine
a0_55|NA|hydroxychlorocquine
a0_55|NA|hydoroxychloroquine
a0_55|NA|hydroxychlororquine
a0_55|NA|hydorxychloroquine
a0_55|NA|hydroxychlroroquine
a0_55|NA|hydroxychlorquine
a0_55|NA|hydrosxychloroquine
a0_55|NA|hydroxychlorooquine
a0_55|NA|hydroxychlorolquine
a0_55|NA|hydroxychlooquine
a0_55|NA|hydrochloroquine
a0_57|NA|COVID 19 respiratory
a0_57|NA|COVID 19 with respiratory
a0_57|NA|COVID 19 w/ respiratory
a0_57|NA|COVID19 respiratory
a0_57|NA|COVID19 with respiratory
a0_57|NA|COVID19 w/ respiratory
a0_57|NA|coronavirus respiratory
a0_57|NA|coronavirus with respiratory
a0_57|NA|coronavirus w/ respiratory
a0_58|NA|COVID19 screening
a0_58|NA|COVID19 screens
a0_58|NA|COVID19 screen
a0_58|NA|screening for COVID19
a0_58|NA|screened for COVID19
a0_58|NA|screens for COVID19
a0_58|NA|screen for COVID19
a0_58|NA|COVID-19 screening
a0_58|NA|COVID-19 screens
a0_58|NA|COVID-19 screen
a0_58|NA|screening for COVID-19
a0_58|NA|screened for COVID-19
a0_58|NA|screens for COVID-19
a0_58|NA|screen for COVID-19
a0_58|NA|COVID screening
a0_58|NA|COVID screens
a0_58|NA|COVID screen
a0_58|NA|screening for COVID
a0_58|NA|screened for COVID
a0_58|NA|screens for COVID
a0_58|NA|screen for COVID
a0_58|NA|novel coronavirus screening
a0_58|NA|novel coronavirus screens
a0_58|NA|novel coronavirus screen
a0_58|NA|screening for novel coronavirus
a0_58|NA|screened for novel coronavirus
a0_58|NA|screens for novel coronavirus
a0_58|NA|screen for novel coronavirus
a0_58|NA|screening for the novel coronavirus
a0_58|NA|screened for the novel coronavirus
a0_58|NA|screens for the novel coronavirus
a0_58|NA|screen for the novel coronavirus
a0_58|NA|coronavirus screening
a0_58|NA|coronavirus screens
a0_58|NA|coronavirus screen
a0_58|NA|screening for coronavirus
a0_58|NA|screened for coronavirus
a0_58|NA|screens for coronavirus
a0_58|NA|screen for coronavirus
a0_58|NA|screening for the coronavirus
a0_58|NA|screened for the coronavirus
a0_58|NA|screens for the coronavirus
a0_58|NA|screen for the coronavirus
a0_59|NA|healthy immune response
a0_59|NA|healthy immune responses
a0_59|NA|normal immune response
a0_59|NA|normal immune responses
a0_59|NA|appropriate immune response
a0_59|NA|appropriate immune responses
a0_59|NA|good immune response
a0_59|NA|good immune responses
a0_59|NA|adequate immune response
a0_59|NA|adequate immune responses
a0_59|NA|healthy immune reaction
a0_59|NA|healthy immune reactions
a0_59|NA|normal immune reaction
a0_59|NA|normal immune reactions
a0_59|NA|appropriate immune reaction
a0_59|NA|appropriate immune reactions
a0_59|NA|good immune reaction
a0_59|NA|good immune reactions
a0_59|NA|adequate immune reaction
a0_59|NA|adequate immune reactions
a0_60|NA|COVID-19 Ab IgG
a0_60|NA|COVID-19 Ab immunoglobulin G
a0_60|NA|COVID-19 antibody IgG
a0_60|NA|COVID-19 antibody immunoglobulin G
a0_60|NA|COVID-19 Ab
a0_60|NA|COVID-19 Abs
a0_60|NA|COVID-19 antibodies
a0_60|NA|COVID-19 antibody
a0_60|NA|immunoglobulin G COVID-19
a0_60|NA|IgG COVID-19
a0_60|NA|immunoglobulin G to COVID-19
a0_60|NA|IgG to COVID-19
a0_60|NA|antibodies to COVID-19
a0_60|NA|antibody to COVID-19
a0_60|NA|Abs to COVID-19
a0_60|NA|Ab to COVID-19
a0_60|NA|COVID19 Ab IgG
a0_60|NA|COVID19 Ab immunoglobulin G
a0_60|NA|COVID19 antibody IgG
a0_60|NA|COVID19 antibody immunoglobulin G
a0_60|NA|COVID19 Ab
a0_60|NA|COVID19 Abs
a0_60|NA|COVID19 antibodies
a0_60|NA|COVID19 antibody
a0_60|NA|immunoglobulin G COVID19
a0_60|NA|IgG COVID19
a0_60|NA|immunoglobulin G to COVID19
a0_60|NA|IgG to COVID19
a0_60|NA|antibodies to COVID19
a0_60|NA|antibody to COVID19
a0_60|NA|Abs to COVID19
a0_60|NA|Ab to COVID19
a0_60|NA|COVID Ab IgG
a0_60|NA|COVID Ab immunoglobulin G
a0_60|NA|COVID antibody IgG
a0_60|NA|COVID antibody immunoglobulin G
a0_60|NA|COVID Ab
a0_60|NA|COVID Abs
a0_60|NA|COVID antibodies
a0_60|NA|COVID antibody
a0_60|NA|immunoglobulin G COVID
a0_60|NA|IgG COVID
a0_60|NA|immunoglobulin G to COVID
a0_60|NA|IgG to COVID
a0_60|NA|antibodies to COVID
a0_60|NA|antibody to COVID
a0_60|NA|Abs to COVID
a0_60|NA|Ab to COVID
a0_60|NA|coronavirus Ab IgG
a0_60|NA|coronavirus Ab immunoglobulin G
a0_60|NA|coronavirus antibody IgG
a0_60|NA|coronavirus antibody immunoglobulin G
a0_60|NA|coronavirus Ab
a0_60|NA|coronavirus Abs
a0_60|NA|coronavirus antibodies
a0_60|NA|coronavirus antibody
a0_60|NA|immunoglobulin G coronavirus
a0_60|NA|IgG coronavirus
a0_60|NA|immunoglobulin G to coronavirus
a0_60|NA|IgG to coronavirus
a0_60|NA|antibodies to coronavirus
a0_60|NA|antibody to coronavirus
a0_60|NA|Abs to coronavirus
a0_60|NA|Ab to coronavirus
a0_60|NA|immunoglobulin G to the coronavirus
a0_60|NA|IgG to the coronavirus
a0_60|NA|antibodies to the coronavirus
a0_60|NA|antibody to the coronavirus
a0_60|NA|Abs to the coronavirus
a0_60|NA|Ab to the coronavirus
a0_60|NA|immunoglobulin G to the novel coronavirus
a0_60|NA|IgG to the novel coronavirus
a0_60|NA|antibodies to the novel coronavirus
a0_60|NA|antibody to the novel coronavirus
a0_60|NA|Abs to the novel coronavirus
a0_60|NA|Ab to the novel coronavirus
a0_61|NA|COVID19 exposure
a0_61|NA|COVID19 exposures
a0_61|NA|exposures to COVID19
a0_61|NA|exposure to COVID19
a0_61|NA|exposing to COVID19
a0_61|NA|exposed to COVID19
a0_61|NA|exposes to COVID19
a0_61|NA|expose to COVID19
a0_61|NA|COVID-19 exposure
a0_61|NA|COVID-19 exposures
a0_61|NA|exposures to COVID-19
a0_61|NA|exposure to COVID-19
a0_61|NA|exposing to COVID-19
a0_61|NA|exposed to COVID-19
a0_61|NA|exposes to COVID-19
a0_61|NA|expose to COVID-19
a0_61|NA|COVID exposure
a0_61|NA|COVID exposures
a0_61|NA|exposures to COVID
a0_61|NA|exposure to COVID
a0_61|NA|exposing to COVID
a0_61|NA|exposed to COVID
a0_61|NA|exposes to COVID
a0_61|NA|expose to COVID
a0_61|NA|novel coronavirus exposure
a0_61|NA|novel coronavirus exposures
a0_61|NA|exposures to the novel coronavirus
a0_61|NA|exposure to the novel coronavirus
a0_61|NA|exposing to the novel coronavirus
a0_61|NA|exposed to the novel coronavirus
a0_61|NA|exposes to the novel coronavirus
a0_61|NA|expose to the novel coronavirus
a0_61|NA|coronavirus exposure
a0_61|NA|coronavirus exposures
a0_61|NA|exposures to the coronavirus
a0_61|NA|exposure to the coronavirus
a0_61|NA|exposing to the coronavirus
a0_61|NA|exposed to the coronavirus
a0_61|NA|exposes to the coronavirus
a0_61|NA|expose to the coronavirus
a0_62|NA|2019 novel coronavirus RNA
a0_62|NA|2019 coronavirus RNA
a0_62|NA|coronavirus RNA
a0_62|NA|COVID-19 RNA
a0_62|NA|COVID19 RNA
a0_62|NA|COVID RNA
a0_63|NA|COVID19 convalescent plasma
a0_63|NA|COVID19 convalescent plasmas
a0_63|NA|COVID19 convalescent serum
a0_63|NA|COVID19 convalescent sera
a0_63|NA|COVID19 convalescent antibodies
a0_63|NA|COVID19 convalescent antibody
a0_63|NA|COVID19 convalescent Abs
a0_63|NA|COVID19 convalescent Ab
a0_63|NA|convalescent COVID19 plasma
a0_63|NA|convalescent COVID19 plasmas
a0_63|NA|convalescent COVID19 serum
a0_63|NA|convalescent COVID19 sera
a0_63|NA|convalescent COVID19 antibodies
a0_63|NA|convalescent COVID19 antibody
a0_63|NA|convalescent COVID19 Abs
a0_63|NA|convalescent COVID19 Ab
a0_63|NA|plasma from recovered COVID19 patients
a0_63|NA|plasma from recovered COVID19 patient
a0_63|NA|plasma from a recovered COVID19 patient
a0_63|NA|serum from recovered COVID19 patients
a0_63|NA|serum from recovered COVID19 patient
a0_63|NA|serum from a recovered COVID19 patient
a0_63|NA|antibodies from recovered COVID19 patients
a0_63|NA|antibodies from recovered COVID19 patient
a0_63|NA|antibodies from a recovered COVID19 patient
a0_63|NA|antibody from recovered COVID19 patients
a0_63|NA|antibody from recovered COVID19 patient
a0_63|NA|antibody from a recovered COVID19 patient
a0_63|NA|Abs from recovered COVID19 patients
a0_63|NA|Abs from recovered COVID19 patient
a0_63|NA|Abs from a recovered COVID19 patient
a0_63|NA|Ab from recovered COVID19 patients
a0_63|NA|Ab from recovered COVID19 patient
a0_63|NA|Ab from a recovered COVID19 patient
a0_65|NA|COVID-19 swab
a0_65|NA|COVID-19 swabbing
a0_65|NA|COVID-19 swabs
a0_65|NA|swabbing for COVID-19
a0_65|NA|swabbed for COVID-19
a0_65|NA|swabs for COVID-19
a0_65|NA|swab for COVID-19
a0_65|NA|swabbing COVID-19
a0_65|NA|swabbed COVID-19
a0_65|NA|swabs COVID-19
a0_65|NA|swab COVID-19
a0_65|NA|COVID19 swab
a0_65|NA|COVID19 swabbed
a0_65|NA|COVID19 swabbing
a0_65|NA|COVID19 swabs
a0_65|NA|swabbing for COVID19
a0_65|NA|swabbed for COVID19
a0_65|NA|swabs for COVID19
a0_65|NA|swab for COVID19
a0_65|NA|swabbing COVID19
a0_65|NA|swabbed COVID19
a0_65|NA|swabs COVID19
a0_65|NA|swab COVID19
a0_65|NA|COVID swab
a0_65|NA|COVID swabbing
a0_65|NA|COVID swabs
a0_65|NA|swabbing for COVID
a0_65|NA|swabbed for COVID
a0_65|NA|swabs for COVID
a0_65|NA|swab for COVID
a0_65|NA|swabbing COVID
a0_65|NA|swabbed COVID
a0_65|NA|swabs COVID
a0_65|NA|swab COVID
a0_65|NA|coronavirus swab
a0_65|NA|coronavirus swabbing
a0_65|NA|coronavirus swabs
a0_65|NA|swabbing for coronavirus
a0_65|NA|swabbed for coronavirus
a0_65|NA|swabs for coronavirus
a0_65|NA|swab for coronavirus
a0_65|NA|swabbing coronavirus
a0_65|NA|swabbed coronavirus
a0_65|NA|swab coronavirus
a0_65|NA|swabs coronavirus
a0_65|NA|novel coronavirus swab
a0_65|NA|novel coronavirus swabbing
a0_65|NA|novel coronavirus swabs
a0_65|NA|swabbing for novel coronavirus
a0_65|NA|swabbed for novel coronavirus
a0_65|NA|swabs for novel coronavirus
a0_65|NA|swab for novel coronavirus
a0_65|NA|swabbing novel coronavirus
a0_65|NA|swabbed novel coronavirus
a0_65|NA|swabs novel coronavirus
a0_65|NA|swab novel coronavirus
a0_65|NA|new coronavirus swab
a0_65|NA|new coronavirus swabbing
a0_65|NA|new coronavirus swabs
a0_65|NA|swabbing for new coronavirus
a0_65|NA|swabbed for new coronavirus
a0_65|NA|swabs for new coronavirus
a0_65|NA|swab for new coronavirus
a0_65|NA|swabbing new coronavirus
a0_65|NA|swabbed new coronavirus
a0_65|NA|swabs new coronavirus
a0_65|NA|swab new coronavirus
a0_65|NA|swabbed for the coronavirus
a0_65|NA|swabbed for the new coronavirus
a0_65|NA|swabbed for the novel coronavirus
a0_65|NA|swabbing for the coronavirus
a0_65|NA|swabbing for the new coronavirus
a0_65|NA|swabbing for the novel coronavirus
a0_65|NA|swabs for the coronavirus
a0_65|NA|swab for the coronavirus
a0_65|NA|swabs for the new coronavirus
a0_65|NA|swab for the new coronavirus
a0_65|NA|swabs for the novel coronavirus
a0_65|NA|swab for the novel coronavirus
a0_66|NA|asymptomatic COVID-19 test positive
a0_66|NA|asymptomatic COVID-19 positive
a0_66|NA|asymptomatic COVID19 test positive
a0_66|NA|asymptomatic COVID19 positive
a0_66|NA|COVID19 asymptomatic postive
a0_66|NA|COVID-19 asymptomatic postive
a0_66|NA|COVID19 postive asymptomatic
a0_66|NA|COVID-19 postive asymptomatic
a0_67|NA|COVID19 testing was negative
a0_67|NA|COVID19 test was negative
a0_67|NA|COVID-19 testing was negative
a0_67|NA|COVID-19 test was negative
a0_67|NA|COVID19 testing was neg
a0_67|NA|COVID19 test was neg
a0_67|NA|COVID-19 testing was neg
a0_67|NA|COVID-19 test was neg
a0_67|NA|COVID19 testing is negative
a0_67|NA|COVID19 test is negative
a0_67|NA|COVID-19 testing is negative
a0_67|NA|COVID-19 test is negative
a0_67|NA|COVID19 testing is neg
a0_67|NA|COVID19 test is neg
a0_67|NA|COVID-19 testing is neg
a0_67|NA|COVID-19 test is neg
a0_67|NA|tested negative COVID19
a0_67|NA|tested negative COVID-19
a0_67|NA|tested negative for COVID19
a0_67|NA|tested negative for COVID-19
a0_67|NA|tested neg COVID19
a0_67|NA|tested neg COVID-19
a0_67|NA|tested neg for COVID19
a0_67|NA|tested neg for COVID-19
a0_67|NA|tested negative for the coronavirus
a0_67|NA|tested negative for the novel coronavirus
a0_67|NA|tested neg for the coronavirus
a0_67|NA|tested neg for the novel coronavirus
a0_67|NA|COVID19 test negative
a0_67|NA|COVID 19 test negative
a0_67|NA|coronavirus test negative
a0_67|NA|COVID19 test neg
a0_67|NA|COVID 19 test neg
a0_67|NA|coronavirus test neg
a0_67|NA|COVID 19 negative
a0_67|NA|COVID19 negative
a0_67|NA|COVID negative
a0_67|NA|2019 novel coronavirus negative
a0_67|NA|COVID 19 PCR negative for 2019 novel coronavirus
a0_67|NA|PCR negative for 2019 novel coronavirus
a0_67|NA|PCR negative for novel coronavirus
a0_67|NA|PCR negative for COVID 19
a0_67|NA|PCR negative for COVID19
a0_67|NA|PCR negative for COVID
a0_67|NA|negative COVID 19 test result
a0_67|NA|negative COVID 19 result
a0_67|NA|negative COVID19 test result
a0_67|NA|negative COVID19 result
a0_67|NA|negative COVID test result
a0_67|NA|negative COVID result
a0_67|NA|negative for 2019 novel coronavirus
a0_67|NA|negative for novel coronavirus
a0_67|NA|negative for COVID 19
a0_67|NA|negative for COVID19
a0_67|NA|negative for COVID
a0_67|NA|negative for 2019 novel coronavirus RNA
a0_67|NA|negative for novel coronavirus RNA
a0_67|NA|negative for COVID 19 RNA
a0_67|NA|negative for COVID19 RNA
a0_67|NA|negative for COVID RNA
a0_67|NA|real time PCR negative for 2019 novel coronavirus
a0_67|NA|real time PCR negative for novel coronavirus
a0_67|NA|real time PCR negative for coronavirus
a0_67|NA|real time PCR negative for COVID 19
a0_67|NA|real time PCR negative for COVID19
a0_67|NA|real time PCR negative for COVID
a0_67|NA|COVID 19 neg
a0_67|NA|COVID19 neg
a0_67|NA|COVID neg
a0_67|NA|2019 novel coronavirus neg
a0_67|NA|COVID 19 PCR neg for 2019 novel coronavirus
a0_67|NA|PCR neg for 2019 novel coronavirus
a0_67|NA|PCR neg for novel coronavirus
a0_67|NA|PCR neg for COVID 19
a0_67|NA|PCR neg for COVID19
a0_67|NA|PCR neg for COVID
a0_67|NA|neg COVID 19 test result
a0_67|NA|neg COVID 19 result
a0_67|NA|neg COVID19 test result
a0_67|NA|neg COVID19 result
a0_67|NA|neg COVID test result
a0_67|NA|neg COVID result
a0_67|NA|neg for 2019 novel coronavirus
a0_67|NA|neg for novel coronavirus
a0_67|NA|neg for COVID 19
a0_67|NA|neg for COVID19
a0_67|NA|neg for COVID
a0_67|NA|neg for 2019 novel coronavirus RNA
a0_67|NA|neg for novel coronavirus RNA
a0_67|NA|neg for COVID 19 RNA
a0_67|NA|neg for COVID19 RNA
a0_67|NA|neg for COVID RNA
a0_67|NA|real time PCR neg for 2019 novel coronavirus
a0_67|NA|real time PCR neg for novel coronavirus
a0_67|NA|real time PCR neg for coronavirus
a0_67|NA|real time PCR neg for COVID 19
a0_67|NA|real time PCR neg for COVID19
a0_67|NA|real time PCR neg for COVID
a0_68|NA|COVID19 convalescent plasma
a0_68|NA|COVID19 convalescent plasmas
a0_68|NA|COVID19 convalescent serum
a0_68|NA|COVID19 convalescent sera
a0_68|NA|COVID19 convalescent antibodies
a0_68|NA|COVID19 convalescent antibody
a0_68|NA|COVID19 convalescent Abs
a0_68|NA|COVID19 convalescent Ab
a0_68|NA|COVID-19 convalescent plasma
a0_68|NA|COVID-19 convalescent plasmas
a0_68|NA|COVID-19 convalescent serum
a0_68|NA|COVID-19 convalescent sera
a0_68|NA|COVID-19 convalescent antibodies
a0_68|NA|COVID-19 convalescent antibody
a0_68|NA|COVID-19 convalescent Abs
a0_68|NA|COVID-19 convalescent Ab
a0_68|NA|convalescent plasma
a0_68|NA|convalescent plasmas
a0_68|NA|convalescent serum
a0_68|NA|convalescent sera
a0_68|NA|convalescent antibodies
a0_68|NA|convalescent antibody
a0_68|NA|convalescent Abs
a0_68|NA|convalescent Ab
a0_69|NA|coronavirus2019
a0_69|NA|coronavirus 2019
a0_69|NA|coronavirus 19
a0_69|NA|COVID-19
a0_69|NA|COVID19
a0_69|NA|COVID
a0_69|NA|corona virus disease 19
a0_69|NA|corona virus disease 2019
a0_69|NA|corona virus disease
a0_69|NA|coronavirus disease 19
a0_69|NA|coronavirus disease 2019
a0_69|NA|coronavirus disease
a0_69|NA|coronavirus
a0_69|NA|CORVID-19
a0_69|NA|CORVID19
a0_69|NA|CORVID
a0_69|NA|CORVIN-19
a0_69|NA|CORVIN19
a0_69|NA|CORVIN
a0_69|NA|COVIN-19
a0_69|NA|COVIN19
a0_69|NA|COVIN
a0_69|NA|CoronavirusDisease
a0_69|NA|COAVID-19
a0_69|NA|COAVID19
a0_69|NA|COAVID
a0_69|NA|COVD-19
a0_69|NA|COVD19
a0_69|NA|COVD
a0_69|NA|CAVIN-19
a0_69|NA|CAVIN19
a0_69|NA|CAVIN
a0_69|NA|novel coronvirus
a0_69|NA|CODIV-19
a0_69|NA|CODIV19
a0_69|NA|CODIV
a0_69|NA|1COVID19
a0_70|NA|COVID-19 signs
a0_70|NA|COVID-19 sign
a0_70|NA|signs of COVID-19
a0_70|NA|sign of COVID-19
a0_70|NA|COVID19 signs
a0_70|NA|COVID19 sign
a0_70|NA|signs of COVID19
a0_70|NA|sign of COVID19
a0_70|NA|COVID signs
a0_70|NA|COVID sign
a0_70|NA|signs of COVID
a0_70|NA|sign of COVID
a0_70|NA|coronavirus signs
a0_70|NA|coronavirus sign
a0_70|NA|signs of coronavirus
a0_70|NA|sign of coronavirus
a0_70|NA|signs of the coronavirus
a0_70|NA|sign of the coronavirus
a0_70|NA|novel signs
a0_70|NA|novel sign
a0_70|NA|signs of novel
a0_70|NA|sign of novel
a0_70|NA|signs of the novel
a0_70|NA|sign of the novel
a0_71|NA|first human vaccine trial
a0_71|NA|first human vaccine trials
a0_71|NA|human vaccine trial
a0_71|NA|human vaccine trials
a0_71|NA|first vaccine trial in humans
a0_71|NA|first vaccine trials in humans
a0_71|NA|vaccine trial in humans
a0_71|NA|vaccine trials in humans
a0_71|NA|vaccine trial
a0_71|NA|vaccine trials
a0_72|NA|coronavirus disease 2019
a0_72|NA|coronavirus disease 19
a0_72|NA|acoronavirus disease
a0_72|NA|COVID-19 disease
a0_72|NA|COVID19 disease
a0_72|NA|COVID disease
a0_72|NA|nCoV-2019
a0_72|NA|nCoV-19
a0_72|NA|nCoV19
a0_72|NA|19-nCoV
a0_72|NA|COVID-19 novel
a0_72|NA|COVID19 novel
a0_72|NA|COVID novel
a0_72|NA|coronavirus COVID-19
a0_72|NA|coronavirus COVID-2019
a0_72|NA|coronavirus COVID19
a0_72|NA|coronavirus COVID2019
a0_72|NA|coronavirus COVID
a0_72|NA|COVID-19 coronavirus
a0_72|NA|COVID19 coronavirus
a0_72|NA|COVID-2019 coronavirus
a0_72|NA|COVID2019 coronavirus
a0_72|NA|COVID coronavirus
a0_72|NA|COVID-19 virus
a0_72|NA|COVID19 virus
a0_72|NA|COVID-2019 virus
a0_72|NA|COVID2019 virus
a0_72|NA|COVID virus
a0_72|NA|SARSCoV-2
a0_72|NA|SARSCoV2
a0_72|NA|SARSCoV
a0_72|NA|novel coronavirus (COVID-19)
a0_72|NA|novel coronavirus (COVID19)
a0_72|NA|novel coronavirus (COVID)
a0_72|NA|novel coronavirus 2019
a0_72|NA|novel coronavirus
a0_72|NA|novel 2019 coronavirus
a0_72|NA|novel 2019 CoV
a0_72|NA|new coronavirus
a0_72|NA|new 2019 coronavirus
a0_72|NA|new 2019 CoV
a0_72|NA|2019 novel coronavirus acute respiratory disease
a0_72|NA|2019 novel coronavirus
a0_72|NA|2019 novel CoV
a0_72|NA|2019 coronavirus acute respiratory disease
a0_72|NA|2019-nCoV acute respiratory disease
a0_72|NA|19 novel coronavirus acute respiratory disease
a0_72|NA|19 novel coronavirus
a0_72|NA|19 novel CoV
a0_72|NA|19 coronavirus acute respiratory disease
a0_72|NA|19-nCoV acute respiratory disease
a0_72|NA|nCoV acute respiratory disease
a0_72|NA|SARS-CoV-2
a0_72|NA|SARS-CoV2
a0_72|NA|SARS-CoV
a0_72|NA|SARS-CoV-19
a0_72|NA|SARS-CoV-2019
a0_72|NA|2019 coronavirus-2
a0_72|NA|2019 coronavirus
a0_72|NA|19 coronavirus-2
a0_72|NA|19 coronavirus
a0_72|NA|severe acute respiratory syndrome coronavirus 2
a0_72|NA|severe acute respiratory syndrome coronavirus
a0_72|NA|SARS-coronavirus 2
a0_72|NA|SARS-coronavirus
a0_72|NA|Corona Virus Disease 19
a0_72|NA|Corona Virus Disease 2019
a0_72|NA|COVID-19 infections
a0_72|NA|COVID19 infections
a0_72|NA|COVID-19 infection
a0_72|NA|COVID19 infection
a0_72|NA|COVID-19
a0_72|NA|COVID19
a0_72|NA|CV19
a0_72|NA|CV-19
a0_72|NA|COVID-2019 infections
a0_72|NA|COVID2019 infections
a0_72|NA|COVID-2019 infection
a0_72|NA|COVID2019 infection
a0_72|NA|COVID-2019
a0_72|NA|CV2019
a0_72|NA|CV-2019
a0_72|NA|2019-nCoV
a0_72|NA|Wuhan coronavirus
a0_72|NA|Wuhan virus
a0_72|NA|coronavirus
a0_72|NA|corona-virus
a0_72|NA|Chinese virus
a0_72|NA|Chinese coronavirus
a0_72|NA|COVID2019
a0_72|NA|corona 2019
a0_72|NA|novel corona
a0_72|NA|U07.1
a0_72|NA|U 07.1
a0_73|NA|coronaviral
a0_73|NA|coronavirus diseases
a0_73|NA|coronavirus disease
a0_73|NA|Coronaviridae
a0_73|NA|coronaviruses
a0_73|NA|coronavirus
a0_73|NA|corona virus diseases
a0_73|NA|corona virus disease
a0_73|NA|Corona viridae
a0_73|NA|corona viruses
a0_73|NA|corona virus
a0_73|NA|CoV
a0_73|NA|CoVs
a0_73|NA|coronoviruses
a0_73|NA|coronovirus
a0_73|NA|coro navirus
a0_73|NA|coronaviruse
a0_73|NA|cornavirus
a0_73|NA|Coronavirinae
a0_73|NA|conronavirus
a0_73|NA|coroanvirus
a0_73|NA|coronvirus
a0_73|NA|coronviruses
a0_73|NA|caronavirus
a0_73|NA|cornoavirus
a0_73|NA|coronoavirus
a0_73|NA|coronaviurs
a0_73|NA|coronaivrus
a0_73|NA|coronavorus
a0_73|NA|coronarvirus
a0_73|NA|coronavirdae
a0_73|NA|coronaviruas
a0_73|NA|coranavirus
a0_73|NA|coronaviru
a0_73|NA|coronavirs
a0_74|NA|shelter in place
a0_74|NA|sheltered in place
a0_74|NA|shelters in place
a0_74|NA|sheltering in place
a0_74|NA|staying at home
a0_74|NA|stays at home
a0_74|NA|stay at home
a0_74|NA|stayed at home
a0_74|NA|staying home
a0_74|NA|stays home
a0_74|NA|stay home
a0_74|NA|stayed home
a0_74|NA|did not leave her home
a0_74|NA|did not leave his home
a0_74|NA|did not leave the home
a0_74|NA|did not leave home
a0_74|NA|did not leave her apartment
a0_74|NA|did not leave his apartment
a0_74|NA|did not leave the apartment
a0_74|NA|did not leave apartment
a0_74|NA|did not leave her house
a0_74|NA|did not leave his house
a0_74|NA|did not leave the house
a0_74|NA|did not leave house
a0_74|NA|did not leave her condo
a0_74|NA|did not leave his condo
a0_74|NA|did not leave the condo
a0_74|NA|did not leave condo
a0_74|NA|didn't leave her apartment
a0_74|NA|didn't leave his apartment
a0_74|NA|didn't leave the apartment
a0_74|NA|didn't leave apartment
a0_74|NA|didn't leave her house
a0_74|NA|didn't leave his house
a0_74|NA|didn't leave the house
a0_74|NA|didn't leave house
a0_74|NA|didn't leave her condo
a0_74|NA|didn't leave his condo
a0_74|NA|didn't leave the condo
a0_74|NA|didn't leave condo
a0_74|NA|not leaving her home
a0_74|NA|not leaving his home
a0_74|NA|not leaving the home
a0_74|NA|not leaving home
a0_74|NA|not leaving her apartment
a0_74|NA|not leaving his apartment
a0_74|NA|not leaving the apartment
a0_74|NA|not leaving apartment
a0_74|NA|not leaving her house
a0_74|NA|not leaving his house
a0_74|NA|not leaving the house
a0_74|NA|not leaving house
a0_74|NA|not leaving her condo
a0_74|NA|not leaving his condo
a0_74|NA|not leaving the condo
a0_74|NA|not leaving condo
a0_75|NA|viral replication
a0_75|NA|viral replications
a0_75|NA|virus replication
a0_75|NA|virus replications
a0_75|NA|replication of viruses
a0_75|NA|replication of virus
a0_75|NA|replication of viral
a0_75|NA|replication of the viruses
a0_75|NA|replication of the virus
a0_75|NA|replication of the viral
a0_75|NA|replicating viruses
a0_75|NA|replicating virus
a0_75|NA|virus replicating
a0_75|NA|virus replicated
a0_75|NA|virus replicates
a0_75|NA|virus replicate
a0_76|NA|incubation period
a0_76|NA|incubation periods
a0_76|NA|incubation time period
a0_76|NA|incubation time periods
a0_76|NA|incubation times
a0_76|NA|incubation time
a0_77|NA|center for a COVID-19 test
a0_77|NA|center for a drive-thru COVID-19 test
a0_77|NA|center for COVID-19 test
a0_77|NA|center for COVID-19 testing
a0_77|NA|center for COVID-19 tests
a0_77|NA|center for drive-thru COVID-19 test
a0_77|NA|center for drive-thru COVID-19 testing
a0_77|NA|center for drive-thru COVID-19 tests
a0_77|NA|centers for a COVID-19 test
a0_77|NA|centers for a drive-thru COVID-19 test
a0_77|NA|centers for COVID-19 test
a0_77|NA|centers for COVID-19 testing
a0_77|NA|centers for COVID-19 tests
a0_77|NA|centers for drive-thru COVID-19 test
a0_77|NA|centers for drive-thru COVID-19 testing
a0_77|NA|centers for drive-thru COVID-19 tests
a0_77|NA|COVID-19 drive-thru
a0_77|NA|COVID-19 drive-thru center
a0_77|NA|COVID-19 drive-thru centers
a0_77|NA|COVID-19 drive-thru location
a0_77|NA|COVID-19 drive-thru locations
a0_77|NA|COVID-19 drive-thru site
a0_77|NA|COVID-19 drive-thru sites
a0_77|NA|COVID-19 drive-thru test
a0_77|NA|COVID-19 drive-thru test center
a0_77|NA|COVID-19 drive-thru test centers
a0_77|NA|COVID-19 drive-thru test location
a0_77|NA|COVID-19 drive-thru test locations
a0_77|NA|COVID-19 drive-thru test site
a0_77|NA|COVID-19 drive-thru test sites
a0_77|NA|COVID-19 drive-thru testing
a0_77|NA|COVID-19 drive-thru testing center
a0_77|NA|COVID-19 drive-thru testing centers
a0_77|NA|COVID-19 drive-thru testing location
a0_77|NA|COVID-19 drive-thru testing locations
a0_77|NA|COVID-19 drive-thru testing site
a0_77|NA|COVID-19 drive-thru testing sites
a0_77|NA|COVID-19 drive-thru tests
a0_77|NA|drive-thru center for a COVID-19 test
a0_77|NA|drive-thru center for COVID-19 test
a0_77|NA|drive-thru center for COVID-19 testing
a0_77|NA|drive-thru center for COVID-19 tests
a0_77|NA|drive-thru centers for a COVID-19 test
a0_77|NA|drive-thru centers for COVID-19 test
a0_77|NA|drive-thru centers for COVID-19 testing
a0_77|NA|drive-thru centers for COVID-19 tests
a0_77|NA|drive-thru location for a COVID-19 test
a0_77|NA|drive-thru location for COVID-19 test
a0_77|NA|drive-thru location for COVID-19 testing
a0_77|NA|drive-thru location for COVID-19 tests
a0_77|NA|drive-thru locations for a COVID-19 test
a0_77|NA|drive-thru locations for COVID-19 test
a0_77|NA|drive-thru locations for COVID-19 testing
a0_77|NA|drive-thru locations for COVID-19 tests
a0_77|NA|drive-thru site for a COVID-19 test
a0_77|NA|drive-thru site for COVID-19 test
a0_77|NA|drive-thru site for COVID-19 testing
a0_77|NA|drive-thru site for COVID-19 tests
a0_77|NA|drive-thru sites for a COVID-19 test
a0_77|NA|drive-thru sites for COVID-19 test
a0_77|NA|drive-thru sites for COVID-19 testing
a0_77|NA|drive-thru sites for COVID-19 tests
a0_77|NA|drive-thru test center for COVID-19
a0_77|NA|drive-thru test centers for COVID-19
a0_77|NA|drive-thru test for COVID-19
a0_77|NA|drive-thru test location for COVID-19
a0_77|NA|drive-thru test locations for COVID-19
a0_77|NA|drive-thru test site for COVID-19
a0_77|NA|drive-thru test sites for COVID-19
a0_77|NA|drive-thru tested for COVID-19
a0_77|NA|drive-thru testing center for COVID-19
a0_77|NA|drive-thru testing centers for COVID-19
a0_77|NA|drive-thru testing for COVID-19
a0_77|NA|drive-thru testing location for COVID-19
a0_77|NA|drive-thru testing locations for COVID-19
a0_77|NA|drive-thru testing site for COVID-19
a0_77|NA|drive-thru testing sites for COVID-19
a0_77|NA|drive-thru tests for COVID-19
a0_77|NA|location for a COVID-19 test
a0_77|NA|location for a drive-thru COVID-19 test
a0_77|NA|location for COVID-19 test
a0_77|NA|location for COVID-19 testing
a0_77|NA|location for COVID-19 tests
a0_77|NA|location for drive-thru COVID-19 test
a0_77|NA|location for drive-thru COVID-19 testing
a0_77|NA|location for drive-thru COVID-19 tests
a0_77|NA|locations for a COVID-19 test
a0_77|NA|locations for a drive-thru COVID-19 test
a0_77|NA|locations for COVID-19 test
a0_77|NA|locations for COVID-19 testing
a0_77|NA|locations for COVID-19 tests
a0_77|NA|locations for drive-thru COVID-19 test
a0_77|NA|locations for drive-thru COVID-19 testing
a0_77|NA|locations for drive-thru COVID-19 tests
a0_77|NA|site for a COVID-19 test
a0_77|NA|site for a drive-thru COVID-19 test
a0_77|NA|site for COVID-19 test
a0_77|NA|site for COVID-19 testing
a0_77|NA|site for COVID-19 tests
a0_77|NA|site for drive-thru COVID-19 test
a0_77|NA|site for drive-thru COVID-19 testing
a0_77|NA|site for drive-thru COVID-19 tests
a0_77|NA|sites for a COVID-19 test
a0_77|NA|sites for a drive-thru COVID-19 test
a0_77|NA|sites for COVID-19 test
a0_77|NA|sites for COVID-19 testing
a0_77|NA|sites for COVID-19 tests
a0_77|NA|sites for drive-thru COVID-19 test
a0_77|NA|sites for drive-thru COVID-19 testing
a0_77|NA|sites for drive-thru COVID-19 tests
a0_77|NA|test center for COVID-19
a0_77|NA|test centers for COVID-19
a0_77|NA|test for COVID-19
a0_77|NA|test location for COVID-19
a0_77|NA|test locations for COVID-19
a0_77|NA|test site for COVID-19
a0_77|NA|test sites for COVID-19
a0_77|NA|tested for COVID-19
a0_77|NA|testing center for COVID-19
a0_77|NA|testing centers for COVID-19
a0_77|NA|testing for COVID-19
a0_77|NA|testing location for COVID-19
a0_77|NA|testing locations for COVID-19
a0_77|NA|testing site for COVID-19
a0_77|NA|testing sites for COVID-19
a0_77|NA|tests for COVID-19
a0_77|NA|center for a COVID19 test
a0_77|NA|center for a drive-thru COVID19 test
a0_77|NA|center for COVID19 test
a0_77|NA|center for COVID19 testing
a0_77|NA|center for COVID19 tests
a0_77|NA|center for drive-thru COVID19 test
a0_77|NA|center for drive-thru COVID19 testing
a0_77|NA|center for drive-thru COVID19 tests
a0_77|NA|centers for a COVID19 test
a0_77|NA|centers for a drive-thru COVID19 test
a0_77|NA|centers for COVID19 test
a0_77|NA|centers for COVID19 testing
a0_77|NA|centers for COVID19 tests
a0_77|NA|centers for drive-thru COVID19 test
a0_77|NA|centers for drive-thru COVID19 testing
a0_77|NA|centers for drive-thru COVID19 tests
a0_77|NA|COVID19 drive-thru
a0_77|NA|COVID19 drive-thru center
a0_77|NA|COVID19 drive-thru centers
a0_77|NA|COVID19 drive-thru location
a0_77|NA|COVID19 drive-thru locations
a0_77|NA|COVID19 drive-thru site
a0_77|NA|COVID19 drive-thru sites
a0_77|NA|COVID19 drive-thru test
a0_77|NA|COVID19 drive-thru test center
a0_77|NA|COVID19 drive-thru test centers
a0_77|NA|COVID19 drive-thru test location
a0_77|NA|COVID19 drive-thru test locations
a0_77|NA|COVID19 drive-thru test site
a0_77|NA|COVID19 drive-thru test sites
a0_77|NA|COVID19 drive-thru testing
a0_77|NA|COVID19 drive-thru testing center
a0_77|NA|COVID19 drive-thru testing centers
a0_77|NA|COVID19 drive-thru testing location
a0_77|NA|COVID19 drive-thru testing locations
a0_77|NA|COVID19 drive-thru testing site
a0_77|NA|COVID19 drive-thru testing sites
a0_77|NA|COVID19 drive-thru tests
a0_77|NA|drive-thru center for a COVID19 test
a0_77|NA|drive-thru center for COVID19 test
a0_77|NA|drive-thru center for COVID19 testing
a0_77|NA|drive-thru center for COVID19 tests
a0_77|NA|drive-thru centers for a COVID19 test
a0_77|NA|drive-thru centers for COVID19 test
a0_77|NA|drive-thru centers for COVID19 testing
a0_77|NA|drive-thru centers for COVID19 tests
a0_77|NA|drive-thru location for a COVID19 test
a0_77|NA|drive-thru location for COVID19 test
a0_77|NA|drive-thru location for COVID19 testing
a0_77|NA|drive-thru location for COVID19 tests
a0_77|NA|drive-thru locations for a COVID19 test
a0_77|NA|drive-thru locations for COVID19 test
a0_77|NA|drive-thru locations for COVID19 testing
a0_77|NA|drive-thru locations for COVID19 tests
a0_77|NA|drive-thru site for a COVID19 test
a0_77|NA|drive-thru site for COVID19 test
a0_77|NA|drive-thru site for COVID19 testing
a0_77|NA|drive-thru site for COVID19 tests
a0_77|NA|drive-thru sites for a COVID19 test
a0_77|NA|drive-thru sites for COVID19 test
a0_77|NA|drive-thru sites for COVID19 testing
a0_77|NA|drive-thru sites for COVID19 tests
a0_77|NA|drive-thru test center for COVID19
a0_77|NA|drive-thru test centers for COVID19
a0_77|NA|drive-thru test for COVID19
a0_77|NA|drive-thru test location for COVID19
a0_77|NA|drive-thru test locations for COVID19
a0_77|NA|drive-thru test site for COVID19
a0_77|NA|drive-thru test sites for COVID19
a0_77|NA|drive-thru tested for COVID19
a0_77|NA|drive-thru testing center for COVID19
a0_77|NA|drive-thru testing centers for COVID19
a0_77|NA|drive-thru testing for COVID19
a0_77|NA|drive-thru testing location for COVID19
a0_77|NA|drive-thru testing locations for COVID19
a0_77|NA|drive-thru testing site for COVID19
a0_77|NA|drive-thru testing sites for COVID19
a0_77|NA|drive-thru tests for COVID19
a0_77|NA|location for a COVID19 test
a0_77|NA|location for a drive-thru COVID19 test
a0_77|NA|location for COVID19 test
a0_77|NA|location for COVID19 testing
a0_77|NA|location for COVID19 tests
a0_77|NA|location for drive-thru COVID19 test
a0_77|NA|location for drive-thru COVID19 testing
a0_77|NA|location for drive-thru COVID19 tests
a0_77|NA|locations for a COVID19 test
a0_77|NA|locations for a drive-thru COVID19 test
a0_77|NA|locations for COVID19 test
a0_77|NA|locations for COVID19 testing
a0_77|NA|locations for COVID19 tests
a0_77|NA|locations for drive-thru COVID19 test
a0_77|NA|locations for drive-thru COVID19 testing
a0_77|NA|locations for drive-thru COVID19 tests
a0_77|NA|site for a COVID19 test
a0_77|NA|site for a drive-thru COVID19 test
a0_77|NA|site for COVID19 test
a0_77|NA|site for COVID19 testing
a0_77|NA|site for COVID19 tests
a0_77|NA|site for drive-thru COVID19 test
a0_77|NA|site for drive-thru COVID19 testing
a0_77|NA|site for drive-thru COVID19 tests
a0_77|NA|sites for a COVID19 test
a0_77|NA|sites for a drive-thru COVID19 test
a0_77|NA|sites for COVID19 test
a0_77|NA|sites for COVID19 testing
a0_77|NA|sites for COVID19 tests
a0_77|NA|sites for drive-thru COVID19 test
a0_77|NA|sites for drive-thru COVID19 testing
a0_77|NA|sites for drive-thru COVID19 tests
a0_77|NA|test center for COVID19
a0_77|NA|test centers for COVID19
a0_77|NA|test for COVID19
a0_77|NA|test location for COVID19
a0_77|NA|test locations for COVID19
a0_77|NA|test site for COVID19
a0_77|NA|test sites for COVID19
a0_77|NA|tested for COVID19
a0_77|NA|testing center for COVID19
a0_77|NA|testing centers for COVID19
a0_77|NA|testing for COVID19
a0_77|NA|testing location for COVID19
a0_77|NA|testing locations for COVID19
a0_77|NA|testing site for COVID19
a0_77|NA|testing sites for COVID19
a0_77|NA|tests for COVID19
a0_77|NA|center for a coronavirus test
a0_77|NA|center for a drive-thru coronavirus test
a0_77|NA|center for coronavirus test
a0_77|NA|center for coronavirus testing
a0_77|NA|center for coronavirus tests
a0_77|NA|center for drive-thru coronavirus test
a0_77|NA|center for drive-thru coronavirus testing
a0_77|NA|center for drive-thru coronavirus tests
a0_77|NA|centers for a coronavirus test
a0_77|NA|centers for a drive-thru coronavirus test
a0_77|NA|centers for coronavirus test
a0_77|NA|centers for coronavirus testing
a0_77|NA|centers for coronavirus tests
a0_77|NA|centers for drive-thru coronavirus test
a0_77|NA|centers for drive-thru coronavirus testing
a0_77|NA|centers for drive-thru coronavirus tests
a0_77|NA|coronavirus drive-thru
a0_77|NA|coronavirus drive-thru center
a0_77|NA|coronavirus drive-thru centers
a0_77|NA|coronavirus drive-thru location
a0_77|NA|coronavirus drive-thru locations
a0_77|NA|coronavirus drive-thru site
a0_77|NA|coronavirus drive-thru sites
a0_77|NA|coronavirus drive-thru test
a0_77|NA|coronavirus drive-thru test center
a0_77|NA|coronavirus drive-thru test centers
a0_77|NA|coronavirus drive-thru test location
a0_77|NA|coronavirus drive-thru test locations
a0_77|NA|coronavirus drive-thru test site
a0_77|NA|coronavirus drive-thru test sites
a0_77|NA|coronavirus drive-thru testing
a0_77|NA|coronavirus drive-thru testing center
a0_77|NA|coronavirus drive-thru testing centers
a0_77|NA|coronavirus drive-thru testing location
a0_77|NA|coronavirus drive-thru testing locations
a0_77|NA|coronavirus drive-thru testing site
a0_77|NA|coronavirus drive-thru testing sites
a0_77|NA|coronavirus drive-thru tests
a0_77|NA|drive-thru center for a coronavirus test
a0_77|NA|drive-thru center for coronavirus test
a0_77|NA|drive-thru center for coronavirus testing
a0_77|NA|drive-thru center for coronavirus tests
a0_77|NA|drive-thru centers for a coronavirus test
a0_77|NA|drive-thru centers for coronavirus test
a0_77|NA|drive-thru centers for coronavirus testing
a0_77|NA|drive-thru centers for coronavirus tests
a0_77|NA|drive-thru location for a coronavirus test
a0_77|NA|drive-thru location for coronavirus test
a0_77|NA|drive-thru location for coronavirus testing
a0_77|NA|drive-thru location for coronavirus tests
a0_77|NA|drive-thru locations for a coronavirus test
a0_77|NA|drive-thru locations for coronavirus test
a0_77|NA|drive-thru locations for coronavirus testing
a0_77|NA|drive-thru locations for coronavirus tests
a0_77|NA|drive-thru site for a coronavirus test
a0_77|NA|drive-thru site for coronavirus test
a0_77|NA|drive-thru site for coronavirus testing
a0_77|NA|drive-thru site for coronavirus tests
a0_77|NA|drive-thru sites for a coronavirus test
a0_77|NA|drive-thru sites for coronavirus test
a0_77|NA|drive-thru sites for coronavirus testing
a0_77|NA|drive-thru sites for coronavirus tests
a0_77|NA|drive-thru test center for coronavirus
a0_77|NA|drive-thru test centers for coronavirus
a0_77|NA|drive-thru test for coronavirus
a0_77|NA|drive-thru test location for coronavirus
a0_77|NA|drive-thru test locations for coronavirus
a0_77|NA|drive-thru test site for coronavirus
a0_77|NA|drive-thru test sites for coronavirus
a0_77|NA|drive-thru tested for coronavirus
a0_77|NA|drive-thru testing center for coronavirus
a0_77|NA|drive-thru testing centers for coronavirus
a0_77|NA|drive-thru testing for coronavirus
a0_77|NA|drive-thru testing location for coronavirus
a0_77|NA|drive-thru testing locations for coronavirus
a0_77|NA|drive-thru testing site for coronavirus
a0_77|NA|drive-thru testing sites for coronavirus
a0_77|NA|drive-thru tests for coronavirus
a0_77|NA|location for a coronavirus test
a0_77|NA|location for a drive-thru coronavirus test
a0_77|NA|location for coronavirus test
a0_77|NA|location for coronavirus testing
a0_77|NA|location for coronavirus tests
a0_77|NA|location for drive-thru coronavirus test
a0_77|NA|location for drive-thru coronavirus testing
a0_77|NA|location for drive-thru coronavirus tests
a0_77|NA|locations for a coronavirus test
a0_77|NA|locations for a drive-thru coronavirus test
a0_77|NA|locations for coronavirus test
a0_77|NA|locations for coronavirus testing
a0_77|NA|locations for coronavirus tests
a0_77|NA|locations for drive-thru coronavirus test
a0_77|NA|locations for drive-thru coronavirus testing
a0_77|NA|locations for drive-thru coronavirus tests
a0_77|NA|site for a coronavirus test
a0_77|NA|site for a drive-thru coronavirus test
a0_77|NA|site for coronavirus test
a0_77|NA|site for coronavirus testing
a0_77|NA|site for coronavirus tests
a0_77|NA|site for drive-thru coronavirus test
a0_77|NA|site for drive-thru coronavirus testing
a0_77|NA|site for drive-thru coronavirus tests
a0_77|NA|sites for a coronavirus test
a0_77|NA|sites for a drive-thru coronavirus test
a0_77|NA|sites for coronavirus test
a0_77|NA|sites for coronavirus testing
a0_77|NA|sites for coronavirus tests
a0_77|NA|sites for drive-thru coronavirus test
a0_77|NA|sites for drive-thru coronavirus testing
a0_77|NA|sites for drive-thru coronavirus tests
a0_77|NA|test center for coronavirus
a0_77|NA|test centers for coronavirus
a0_77|NA|test for coronavirus
a0_77|NA|test location for coronavirus
a0_77|NA|test locations for coronavirus
a0_77|NA|test site for coronavirus
a0_77|NA|test sites for coronavirus
a0_77|NA|tested for coronavirus
a0_77|NA|testing center for coronavirus
a0_77|NA|testing centers for coronavirus
a0_77|NA|testing for coronavirus
a0_77|NA|testing location for coronavirus
a0_77|NA|testing locations for coronavirus
a0_77|NA|testing site for coronavirus
a0_77|NA|testing sites for coronavirus
a0_77|NA|tests for coronavirus
a0_77|NA|center for a drive-through COVID-19 test
a0_77|NA|center for drive-through COVID-19 test
a0_77|NA|center for drive-through COVID-19 testing
a0_77|NA|center for drive-through COVID-19 tests
a0_77|NA|centers for a drive-through COVID-19 test
a0_77|NA|centers for drive-through COVID-19 test
a0_77|NA|centers for drive-through COVID-19 testing
a0_77|NA|centers for drive-through COVID-19 tests
a0_77|NA|COVID-19 drive-through
a0_77|NA|COVID-19 drive-through center
a0_77|NA|COVID-19 drive-through centers
a0_77|NA|COVID-19 drive-through location
a0_77|NA|COVID-19 drive-through locations
a0_77|NA|COVID-19 drive-through site
a0_77|NA|COVID-19 drive-through sites
a0_77|NA|COVID-19 drive-through test
a0_77|NA|COVID-19 drive-through test center
a0_77|NA|COVID-19 drive-through test centers
a0_77|NA|COVID-19 drive-through test location
a0_77|NA|COVID-19 drive-through test locations
a0_77|NA|COVID-19 drive-through test site
a0_77|NA|COVID-19 drive-through test sites
a0_77|NA|COVID-19 drive-through testing
a0_77|NA|COVID-19 drive-through testing center
a0_77|NA|COVID-19 drive-through testing centers
a0_77|NA|COVID-19 drive-through testing location
a0_77|NA|COVID-19 drive-through testing locations
a0_77|NA|COVID-19 drive-through testing site
a0_77|NA|COVID-19 drive-through testing sites
a0_77|NA|COVID-19 drive-through tests
a0_77|NA|drive-through center for a COVID-19 test
a0_77|NA|drive-through center for COVID-19 test
a0_77|NA|drive-through center for COVID-19 testing
a0_77|NA|drive-through center for COVID-19 tests
a0_77|NA|drive-through centers for a COVID-19 test
a0_77|NA|drive-through centers for COVID-19 test
a0_77|NA|drive-through centers for COVID-19 testing
a0_77|NA|drive-through centers for COVID-19 tests
a0_77|NA|drive-through location for a COVID-19 test
a0_77|NA|drive-through location for COVID-19 test
a0_77|NA|drive-through location for COVID-19 testing
a0_77|NA|drive-through location for COVID-19 tests
a0_77|NA|drive-through locations for a COVID-19 test
a0_77|NA|drive-through locations for COVID-19 test
a0_77|NA|drive-through locations for COVID-19 testing
a0_77|NA|drive-through locations for COVID-19 tests
a0_77|NA|drive-through site for a COVID-19 test
a0_77|NA|drive-through site for COVID-19 test
a0_77|NA|drive-through site for COVID-19 testing
a0_77|NA|drive-through site for COVID-19 tests
a0_77|NA|drive-through sites for a COVID-19 test
a0_77|NA|drive-through sites for COVID-19 test
a0_77|NA|drive-through sites for COVID-19 testing
a0_77|NA|drive-through sites for COVID-19 tests
a0_77|NA|drive-through test center for COVID-19
a0_77|NA|drive-through test centers for COVID-19
a0_77|NA|drive-through test for COVID-19
a0_77|NA|drive-through test location for COVID-19
a0_77|NA|drive-through test locations for COVID-19
a0_77|NA|drive-through test site for COVID-19
a0_77|NA|drive-through test sites for COVID-19
a0_77|NA|drive-through tested for COVID-19
a0_77|NA|drive-through testing center for COVID-19
a0_77|NA|drive-through testing centers for COVID-19
a0_77|NA|drive-through testing for COVID-19
a0_77|NA|drive-through testing location for COVID-19
a0_77|NA|drive-through testing locations for COVID-19
a0_77|NA|drive-through testing site for COVID-19
a0_77|NA|drive-through testing sites for COVID-19
a0_77|NA|drive-through tests for COVID-19
a0_77|NA|location for a drive-through COVID-19 test
a0_77|NA|location for drive-through COVID-19 test
a0_77|NA|location for drive-through COVID-19 testing
a0_77|NA|location for drive-through COVID-19 tests
a0_77|NA|locations for a drive-through COVID-19 test
a0_77|NA|locations for drive-through COVID-19 test
a0_77|NA|locations for drive-through COVID-19 testing
a0_77|NA|locations for drive-through COVID-19 tests
a0_77|NA|site for a drive-through COVID-19 test
a0_77|NA|site for drive-through COVID-19 test
a0_77|NA|site for drive-through COVID-19 testing
a0_77|NA|site for drive-through COVID-19 tests
a0_77|NA|sites for a drive-through COVID-19 test
a0_77|NA|sites for drive-through COVID-19 test
a0_77|NA|sites for drive-through COVID-19 testing
a0_77|NA|sites for drive-through COVID-19 tests
a0_77|NA|center for a drive-through COVID19 test
a0_77|NA|center for drive-through COVID19 test
a0_77|NA|center for drive-through COVID19 testing
a0_77|NA|center for drive-through COVID19 tests
a0_77|NA|centers for a drive-through COVID19 test
a0_77|NA|centers for drive-through COVID19 test
a0_77|NA|centers for drive-through COVID19 testing
a0_77|NA|centers for drive-through COVID19 tests
a0_77|NA|COVID19 drive-through
a0_77|NA|COVID19 drive-through center
a0_77|NA|COVID19 drive-through centers
a0_77|NA|COVID19 drive-through location
a0_77|NA|COVID19 drive-through locations
a0_77|NA|COVID19 drive-through site
a0_77|NA|COVID19 drive-through sites
a0_77|NA|COVID19 drive-through test
a0_77|NA|COVID19 drive-through test center
a0_77|NA|COVID19 drive-through test centers
a0_77|NA|COVID19 drive-through test location
a0_77|NA|COVID19 drive-through test locations
a0_77|NA|COVID19 drive-through test site
a0_77|NA|COVID19 drive-through test sites
a0_77|NA|COVID19 drive-through testing
a0_77|NA|COVID19 drive-through testing center
a0_77|NA|COVID19 drive-through testing centers
a0_77|NA|COVID19 drive-through testing location
a0_77|NA|COVID19 drive-through testing locations
a0_77|NA|COVID19 drive-through testing site
a0_77|NA|COVID19 drive-through testing sites
a0_77|NA|COVID19 drive-through tests
a0_77|NA|drive-through center for a COVID19 test
a0_77|NA|drive-through center for COVID19 test
a0_77|NA|drive-through center for COVID19 testing
a0_77|NA|drive-through center for COVID19 tests
a0_77|NA|drive-through centers for a COVID19 test
a0_77|NA|drive-through centers for COVID19 test
a0_77|NA|drive-through centers for COVID19 testing
a0_77|NA|drive-through centers for COVID19 tests
a0_77|NA|drive-through location for a COVID19 test
a0_77|NA|drive-through location for COVID19 test
a0_77|NA|drive-through location for COVID19 testing
a0_77|NA|drive-through location for COVID19 tests
a0_77|NA|drive-through locations for a COVID19 test
a0_77|NA|drive-through locations for COVID19 test
a0_77|NA|drive-through locations for COVID19 testing
a0_77|NA|drive-through locations for COVID19 tests
a0_77|NA|drive-through site for a COVID19 test
a0_77|NA|drive-through site for COVID19 test
a0_77|NA|drive-through site for COVID19 testing
a0_77|NA|drive-through site for COVID19 tests
a0_77|NA|drive-through sites for a COVID19 test
a0_77|NA|drive-through sites for COVID19 test
a0_77|NA|drive-through sites for COVID19 testing
a0_77|NA|drive-through sites for COVID19 tests
a0_77|NA|drive-through test center for COVID19
a0_77|NA|drive-through test centers for COVID19
a0_77|NA|drive-through test for COVID19
a0_77|NA|drive-through test location for COVID19
a0_77|NA|drive-through test locations for COVID19
a0_77|NA|drive-through test site for COVID19
a0_77|NA|drive-through test sites for COVID19
a0_77|NA|drive-through tested for COVID19
a0_77|NA|drive-through testing center for COVID19
a0_77|NA|drive-through testing centers for COVID19
a0_77|NA|drive-through testing for COVID19
a0_77|NA|drive-through testing location for COVID19
a0_77|NA|drive-through testing locations for COVID19
a0_77|NA|drive-through testing site for COVID19
a0_77|NA|drive-through testing sites for COVID19
a0_77|NA|drive-through tests for COVID19
a0_77|NA|location for a drive-through COVID19 test
a0_77|NA|location for drive-through COVID19 test
a0_77|NA|location for drive-through COVID19 testing
a0_77|NA|location for drive-through COVID19 tests
a0_77|NA|locations for a drive-through COVID19 test
a0_77|NA|locations for drive-through COVID19 test
a0_77|NA|locations for drive-through COVID19 testing
a0_77|NA|locations for drive-through COVID19 tests
a0_77|NA|site for a drive-through COVID19 test
a0_77|NA|site for drive-through COVID19 test
a0_77|NA|site for drive-through COVID19 testing
a0_77|NA|site for drive-through COVID19 tests
a0_77|NA|sites for a drive-through COVID19 test
a0_77|NA|sites for drive-through COVID19 test
a0_77|NA|sites for drive-through COVID19 testing
a0_77|NA|sites for drive-through COVID19 tests
a0_77|NA|center for a drive-through coronavirus test
a0_77|NA|center for drive-through coronavirus test
a0_77|NA|center for drive-through coronavirus testing
a0_77|NA|center for drive-through coronavirus tests
a0_77|NA|centers for a drive-through coronavirus test
a0_77|NA|centers for drive-through coronavirus test
a0_77|NA|centers for drive-through coronavirus testing
a0_77|NA|centers for drive-through coronavirus tests
a0_77|NA|coronavirus drive-through
a0_77|NA|coronavirus drive-through center
a0_77|NA|coronavirus drive-through centers
a0_77|NA|coronavirus drive-through location
a0_77|NA|coronavirus drive-through locations
a0_77|NA|coronavirus drive-through site
a0_77|NA|coronavirus drive-through sites
a0_77|NA|coronavirus drive-through test
a0_77|NA|coronavirus drive-through test center
a0_77|NA|coronavirus drive-through test centers
a0_77|NA|coronavirus drive-through test location
a0_77|NA|coronavirus drive-through test locations
a0_77|NA|coronavirus drive-through test site
a0_77|NA|coronavirus drive-through test sites
a0_77|NA|coronavirus drive-through testing
a0_77|NA|coronavirus drive-through testing center
a0_77|NA|coronavirus drive-through testing centers
a0_77|NA|coronavirus drive-through testing location
a0_77|NA|coronavirus drive-through testing locations
a0_77|NA|coronavirus drive-through testing site
a0_77|NA|coronavirus drive-through testing sites
a0_77|NA|coronavirus drive-through tests
a0_77|NA|drive-through center for a coronavirus test
a0_77|NA|drive-through center for coronavirus test
a0_77|NA|drive-through center for coronavirus testing
a0_77|NA|drive-through center for coronavirus tests
a0_77|NA|drive-through centers for a coronavirus test
a0_77|NA|drive-through centers for coronavirus test
a0_77|NA|drive-through centers for coronavirus testing
a0_77|NA|drive-through centers for coronavirus tests
a0_77|NA|drive-through location for a coronavirus test
a0_77|NA|drive-through location for coronavirus test
a0_77|NA|drive-through location for coronavirus testing
a0_77|NA|drive-through location for coronavirus tests
a0_77|NA|drive-through locations for a coronavirus test
a0_77|NA|drive-through locations for coronavirus test
a0_77|NA|drive-through locations for coronavirus testing
a0_77|NA|drive-through locations for coronavirus tests
a0_77|NA|drive-through site for a coronavirus test
a0_77|NA|drive-through site for coronavirus test
a0_77|NA|drive-through site for coronavirus testing
a0_77|NA|drive-through site for coronavirus tests
a0_77|NA|drive-through sites for a coronavirus test
a0_77|NA|drive-through sites for coronavirus test
a0_77|NA|drive-through sites for coronavirus testing
a0_77|NA|drive-through sites for coronavirus tests
a0_77|NA|drive-through test center for coronavirus
a0_77|NA|drive-through test centers for coronavirus
a0_77|NA|drive-through test for coronavirus
a0_77|NA|drive-through test location for coronavirus
a0_77|NA|drive-through test locations for coronavirus
a0_77|NA|drive-through test site for coronavirus
a0_77|NA|drive-through test sites for coronavirus
a0_77|NA|drive-through tested for coronavirus
a0_77|NA|drive-through testing center for coronavirus
a0_77|NA|drive-through testing centers for coronavirus
a0_77|NA|drive-through testing for coronavirus
a0_77|NA|drive-through testing location for coronavirus
a0_77|NA|drive-through testing locations for coronavirus
a0_77|NA|drive-through testing site for coronavirus
a0_77|NA|drive-through testing sites for coronavirus
a0_77|NA|drive-through tests for coronavirus
a0_77|NA|location for a drive-through coronavirus test
a0_77|NA|location for drive-through coronavirus test
a0_77|NA|location for drive-through coronavirus testing
a0_77|NA|location for drive-through coronavirus tests
a0_77|NA|locations for a drive-through coronavirus test
a0_77|NA|locations for drive-through coronavirus test
a0_77|NA|locations for drive-through coronavirus testing
a0_77|NA|locations for drive-through coronavirus tests
a0_77|NA|site for a drive-through coronavirus test
a0_77|NA|site for drive-through coronavirus test
a0_77|NA|site for drive-through coronavirus testing
a0_77|NA|site for drive-through coronavirus tests
a0_77|NA|sites for a drive-through coronavirus test
a0_77|NA|sites for drive-through coronavirus test
a0_77|NA|sites for drive-through coronavirus testing
a0_77|NA|sites for drive-through coronavirus tests
a0_77|NA|center for a drive-by COVID-19 test
a0_77|NA|center for drive-by COVID-19 test
a0_77|NA|center for drive-by COVID-19 testing
a0_77|NA|center for drive-by COVID-19 tests
a0_77|NA|centers for a drive-by COVID-19 test
a0_77|NA|centers for drive-by COVID-19 test
a0_77|NA|centers for drive-by COVID-19 testing
a0_77|NA|centers for drive-by COVID-19 tests
a0_77|NA|COVID-19 drive-by
a0_77|NA|COVID-19 drive-by center
a0_77|NA|COVID-19 drive-by centers
a0_77|NA|COVID-19 drive-by location
a0_77|NA|COVID-19 drive-by locations
a0_77|NA|COVID-19 drive-by site
a0_77|NA|COVID-19 drive-by sites
a0_77|NA|COVID-19 drive-by test
a0_77|NA|COVID-19 drive-by test center
a0_77|NA|COVID-19 drive-by test centers
a0_77|NA|COVID-19 drive-by test location
a0_77|NA|COVID-19 drive-by test locations
a0_77|NA|COVID-19 drive-by test site
a0_77|NA|COVID-19 drive-by test sites
a0_77|NA|COVID-19 drive-by testing
a0_77|NA|COVID-19 drive-by testing center
a0_77|NA|COVID-19 drive-by testing centers
a0_77|NA|COVID-19 drive-by testing location
a0_77|NA|COVID-19 drive-by testing locations
a0_77|NA|COVID-19 drive-by testing site
a0_77|NA|COVID-19 drive-by testing sites
a0_77|NA|COVID-19 drive-by tests
a0_77|NA|drive-by center for a COVID-19 test
a0_77|NA|drive-by center for COVID-19 test
a0_77|NA|drive-by center for COVID-19 testing
a0_77|NA|drive-by center for COVID-19 tests
a0_77|NA|drive-by centers for a COVID-19 test
a0_77|NA|drive-by centers for COVID-19 test
a0_77|NA|drive-by centers for COVID-19 testing
a0_77|NA|drive-by centers for COVID-19 tests
a0_77|NA|drive-by location for a COVID-19 test
a0_77|NA|drive-by location for COVID-19 test
a0_77|NA|drive-by location for COVID-19 testing
a0_77|NA|drive-by location for COVID-19 tests
a0_77|NA|drive-by locations for a COVID-19 test
a0_77|NA|drive-by locations for COVID-19 test
a0_77|NA|drive-by locations for COVID-19 testing
a0_77|NA|drive-by locations for COVID-19 tests
a0_77|NA|drive-by site for a COVID-19 test
a0_77|NA|drive-by site for COVID-19 test
a0_77|NA|drive-by site for COVID-19 testing
a0_77|NA|drive-by site for COVID-19 tests
a0_77|NA|drive-by sites for a COVID-19 test
a0_77|NA|drive-by sites for COVID-19 test
a0_77|NA|drive-by sites for COVID-19 testing
a0_77|NA|drive-by sites for COVID-19 tests
a0_77|NA|drive-by test center for COVID-19
a0_77|NA|drive-by test centers for COVID-19
a0_77|NA|drive-by test for COVID-19
a0_77|NA|drive-by test location for COVID-19
a0_77|NA|drive-by test locations for COVID-19
a0_77|NA|drive-by test site for COVID-19
a0_77|NA|drive-by test sites for COVID-19
a0_77|NA|drive-by tested for COVID-19
a0_77|NA|drive-by testing center for COVID-19
a0_77|NA|drive-by testing centers for COVID-19
a0_77|NA|drive-by testing for COVID-19
a0_77|NA|drive-by testing location for COVID-19
a0_77|NA|drive-by testing locations for COVID-19
a0_77|NA|drive-by testing site for COVID-19
a0_77|NA|drive-by testing sites for COVID-19
a0_77|NA|drive-by tests for COVID-19
a0_77|NA|location for a drive-by COVID-19 test
a0_77|NA|location for drive-by COVID-19 test
a0_77|NA|location for drive-by COVID-19 testing
a0_77|NA|location for drive-by COVID-19 tests
a0_77|NA|locations for a drive-by COVID-19 test
a0_77|NA|locations for drive-by COVID-19 test
a0_77|NA|locations for drive-by COVID-19 testing
a0_77|NA|locations for drive-by COVID-19 tests
a0_77|NA|site for a drive-by COVID-19 test
a0_77|NA|site for drive-by COVID-19 test
a0_77|NA|site for drive-by COVID-19 testing
a0_77|NA|site for drive-by COVID-19 tests
a0_77|NA|sites for a drive-by COVID-19 test
a0_77|NA|sites for drive-by COVID-19 test
a0_77|NA|sites for drive-by COVID-19 testing
a0_77|NA|sites for drive-by COVID-19 tests
a0_77|NA|center for a drive-by COVID19 test
a0_77|NA|center for drive-by COVID19 test
a0_77|NA|center for drive-by COVID19 testing
a0_77|NA|center for drive-by COVID19 tests
a0_77|NA|centers for a drive-by COVID19 test
a0_77|NA|centers for drive-by COVID19 test
a0_77|NA|centers for drive-by COVID19 testing
a0_77|NA|centers for drive-by COVID19 tests
a0_77|NA|COVID19 drive-by
a0_77|NA|COVID19 drive-by center
a0_77|NA|COVID19 drive-by centers
a0_77|NA|COVID19 drive-by location
a0_77|NA|COVID19 drive-by locations
a0_77|NA|COVID19 drive-by site
a0_77|NA|COVID19 drive-by sites
a0_77|NA|COVID19 drive-by test
a0_77|NA|COVID19 drive-by test center
a0_77|NA|COVID19 drive-by test centers
a0_77|NA|COVID19 drive-by test location
a0_77|NA|COVID19 drive-by test locations
a0_77|NA|COVID19 drive-by test site
a0_77|NA|COVID19 drive-by test sites
a0_77|NA|COVID19 drive-by testing
a0_77|NA|COVID19 drive-by testing center
a0_77|NA|COVID19 drive-by testing centers
a0_77|NA|COVID19 drive-by testing location
a0_77|NA|COVID19 drive-by testing locations
a0_77|NA|COVID19 drive-by testing site
a0_77|NA|COVID19 drive-by testing sites
a0_77|NA|COVID19 drive-by tests
a0_77|NA|drive-by center for a COVID19 test
a0_77|NA|drive-by center for COVID19 test
a0_77|NA|drive-by center for COVID19 testing
a0_77|NA|drive-by center for COVID19 tests
a0_77|NA|drive-by centers for a COVID19 test
a0_77|NA|drive-by centers for COVID19 test
a0_77|NA|drive-by centers for COVID19 testing
a0_77|NA|drive-by centers for COVID19 tests
a0_77|NA|drive-by location for a COVID19 test
a0_77|NA|drive-by location for COVID19 test
a0_77|NA|drive-by location for COVID19 testing
a0_77|NA|drive-by location for COVID19 tests
a0_77|NA|drive-by locations for a COVID19 test
a0_77|NA|drive-by locations for COVID19 test
a0_77|NA|drive-by locations for COVID19 testing
a0_77|NA|drive-by locations for COVID19 tests
a0_77|NA|drive-by site for a COVID19 test
a0_77|NA|drive-by site for COVID19 test
a0_77|NA|drive-by site for COVID19 testing
a0_77|NA|drive-by site for COVID19 tests
a0_77|NA|drive-by sites for a COVID19 test
a0_77|NA|drive-by sites for COVID19 test
a0_77|NA|drive-by sites for COVID19 testing
a0_77|NA|drive-by sites for COVID19 tests
a0_77|NA|drive-by test center for COVID19
a0_77|NA|drive-by test centers for COVID19
a0_77|NA|drive-by test for COVID19
a0_77|NA|drive-by test location for COVID19
a0_77|NA|drive-by test locations for COVID19
a0_77|NA|drive-by test site for COVID19
a0_77|NA|drive-by test sites for COVID19
a0_77|NA|drive-by tested for COVID19
a0_77|NA|drive-by testing center for COVID19
a0_77|NA|drive-by testing centers for COVID19
a0_77|NA|drive-by testing for COVID19
a0_77|NA|drive-by testing location for COVID19
a0_77|NA|drive-by testing locations for COVID19
a0_77|NA|drive-by testing site for COVID19
a0_77|NA|drive-by testing sites for COVID19
a0_77|NA|drive-by tests for COVID19
a0_77|NA|location for a drive-by COVID19 test
a0_77|NA|location for drive-by COVID19 test
a0_77|NA|location for drive-by COVID19 testing
a0_77|NA|location for drive-by COVID19 tests
a0_77|NA|locations for a drive-by COVID19 test
a0_77|NA|locations for drive-by COVID19 test
a0_77|NA|locations for drive-by COVID19 testing
a0_77|NA|locations for drive-by COVID19 tests
a0_77|NA|site for a drive-by COVID19 test
a0_77|NA|site for drive-by COVID19 test
a0_77|NA|site for drive-by COVID19 testing
a0_77|NA|site for drive-by COVID19 tests
a0_77|NA|sites for a drive-by COVID19 test
a0_77|NA|sites for drive-by COVID19 test
a0_77|NA|sites for drive-by COVID19 testing
a0_77|NA|sites for drive-by COVID19 tests
a0_77|NA|center for a drive-by coronavirus test
a0_77|NA|center for drive-by coronavirus test
a0_77|NA|center for drive-by coronavirus testing
a0_77|NA|center for drive-by coronavirus tests
a0_77|NA|centers for a drive-by coronavirus test
a0_77|NA|centers for drive-by coronavirus test
a0_77|NA|centers for drive-by coronavirus testing
a0_77|NA|centers for drive-by coronavirus tests
a0_77|NA|coronavirus drive-by
a0_77|NA|coronavirus drive-by center
a0_77|NA|coronavirus drive-by centers
a0_77|NA|coronavirus drive-by location
a0_77|NA|coronavirus drive-by locations
a0_77|NA|coronavirus drive-by site
a0_77|NA|coronavirus drive-by sites
a0_77|NA|coronavirus drive-by test
a0_77|NA|coronavirus drive-by test center
a0_77|NA|coronavirus drive-by test centers
a0_77|NA|coronavirus drive-by test location
a0_77|NA|coronavirus drive-by test locations
a0_77|NA|coronavirus drive-by test site
a0_77|NA|coronavirus drive-by test sites
a0_77|NA|coronavirus drive-by testing
a0_77|NA|coronavirus drive-by testing center
a0_77|NA|coronavirus drive-by testing centers
a0_77|NA|coronavirus drive-by testing location
a0_77|NA|coronavirus drive-by testing locations
a0_77|NA|coronavirus drive-by testing site
a0_77|NA|coronavirus drive-by testing sites
a0_77|NA|coronavirus drive-by tests
a0_77|NA|drive-by center for a coronavirus test
a0_77|NA|drive-by center for coronavirus test
a0_77|NA|drive-by center for coronavirus testing
a0_77|NA|drive-by center for coronavirus tests
a0_77|NA|drive-by centers for a coronavirus test
a0_77|NA|drive-by centers for coronavirus test
a0_77|NA|drive-by centers for coronavirus testing
a0_77|NA|drive-by centers for coronavirus tests
a0_77|NA|drive-by location for a coronavirus test
a0_77|NA|drive-by location for coronavirus test
a0_77|NA|drive-by location for coronavirus testing
a0_77|NA|drive-by location for coronavirus tests
a0_77|NA|drive-by locations for a coronavirus test
a0_77|NA|drive-by locations for coronavirus test
a0_77|NA|drive-by locations for coronavirus testing
a0_77|NA|drive-by locations for coronavirus tests
a0_77|NA|drive-by site for a coronavirus test
a0_77|NA|drive-by site for coronavirus test
a0_77|NA|drive-by site for coronavirus testing
a0_77|NA|drive-by site for coronavirus tests
a0_77|NA|drive-by sites for a coronavirus test
a0_77|NA|drive-by sites for coronavirus test
a0_77|NA|drive-by sites for coronavirus testing
a0_77|NA|drive-by sites for coronavirus tests
a0_77|NA|drive-by test center for coronavirus
a0_77|NA|drive-by test centers for coronavirus
a0_77|NA|drive-by test for coronavirus
a0_77|NA|drive-by test location for coronavirus
a0_77|NA|drive-by test locations for coronavirus
a0_77|NA|drive-by test site for coronavirus
a0_77|NA|drive-by test sites for coronavirus
a0_77|NA|drive-by tested for coronavirus
a0_77|NA|drive-by testing center for coronavirus
a0_77|NA|drive-by testing centers for coronavirus
a0_77|NA|drive-by testing for coronavirus
a0_77|NA|drive-by testing location for coronavirus
a0_77|NA|drive-by testing locations for coronavirus
a0_77|NA|drive-by testing site for coronavirus
a0_77|NA|drive-by testing sites for coronavirus
a0_77|NA|drive-by tests for coronavirus
a0_77|NA|location for a drive-by coronavirus test
a0_77|NA|location for drive-by coronavirus test
a0_77|NA|location for drive-by coronavirus testing
a0_77|NA|location for drive-by coronavirus tests
a0_77|NA|locations for a drive-by coronavirus test
a0_77|NA|locations for drive-by coronavirus test
a0_77|NA|locations for drive-by coronavirus testing
a0_77|NA|locations for drive-by coronavirus tests
a0_77|NA|site for a drive-by coronavirus test
a0_77|NA|site for drive-by coronavirus test
a0_77|NA|site for drive-by coronavirus testing
a0_77|NA|site for drive-by coronavirus tests
a0_77|NA|sites for a drive-by coronavirus test
a0_77|NA|sites for drive-by coronavirus test
a0_77|NA|sites for drive-by coronavirus testing
a0_77|NA|sites for drive-by coronavirus tests
a0_77|NA|center for a COVID test
a0_77|NA|center for a drive-thru COVID test
a0_77|NA|center for COVID test
a0_77|NA|center for COVID testing
a0_77|NA|center for COVID tests
a0_77|NA|center for drive-thru COVID test
a0_77|NA|center for drive-thru COVID testing
a0_77|NA|center for drive-thru COVID tests
a0_77|NA|centers for a COVID test
a0_77|NA|centers for a drive-thru COVID test
a0_77|NA|centers for COVID test
a0_77|NA|centers for COVID testing
a0_77|NA|centers for COVID tests
a0_77|NA|centers for drive-thru COVID test
a0_77|NA|centers for drive-thru COVID testing
a0_77|NA|centers for drive-thru COVID tests
a0_77|NA|COVID drive-thru
a0_77|NA|COVID drive-thru center
a0_77|NA|COVID drive-thru centers
a0_77|NA|COVID drive-thru location
a0_77|NA|COVID drive-thru locations
a0_77|NA|COVID drive-thru site
a0_77|NA|COVID drive-thru sites
a0_77|NA|COVID drive-thru test
a0_77|NA|COVID drive-thru test center
a0_77|NA|COVID drive-thru test centers
a0_77|NA|COVID drive-thru test location
a0_77|NA|COVID drive-thru test locations
a0_77|NA|COVID drive-thru test site
a0_77|NA|COVID drive-thru test sites
a0_77|NA|COVID drive-thru testing
a0_77|NA|COVID drive-thru testing center
a0_77|NA|COVID drive-thru testing centers
a0_77|NA|COVID drive-thru testing location
a0_77|NA|COVID drive-thru testing locations
a0_77|NA|COVID drive-thru testing site
a0_77|NA|COVID drive-thru testing sites
a0_77|NA|COVID drive-thru tests
a0_77|NA|drive-thru center for a COVID test
a0_77|NA|drive-thru center for COVID test
a0_77|NA|drive-thru center for COVID testing
a0_77|NA|drive-thru center for COVID tests
a0_77|NA|drive-thru centers for a COVID test
a0_77|NA|drive-thru centers for COVID test
a0_77|NA|drive-thru centers for COVID testing
a0_77|NA|drive-thru centers for COVID tests
a0_77|NA|drive-thru location for a COVID test
a0_77|NA|drive-thru location for COVID test
a0_77|NA|drive-thru location for COVID testing
a0_77|NA|drive-thru location for COVID tests
a0_77|NA|drive-thru locations for a COVID test
a0_77|NA|drive-thru locations for COVID test
a0_77|NA|drive-thru locations for COVID testing
a0_77|NA|drive-thru locations for COVID tests
a0_77|NA|drive-thru site for a COVID test
a0_77|NA|drive-thru site for COVID test
a0_77|NA|drive-thru site for COVID testing
a0_77|NA|drive-thru site for COVID tests
a0_77|NA|drive-thru sites for a COVID test
a0_77|NA|drive-thru sites for COVID test
a0_77|NA|drive-thru sites for COVID testing
a0_77|NA|drive-thru sites for COVID tests
a0_77|NA|drive-thru test center for COVID
a0_77|NA|drive-thru test centers for COVID
a0_77|NA|drive-thru test for COVID
a0_77|NA|drive-thru test location for COVID
a0_77|NA|drive-thru test locations for COVID
a0_77|NA|drive-thru test site for COVID
a0_77|NA|drive-thru test sites for COVID
a0_77|NA|drive-thru tested for COVID
a0_77|NA|drive-thru testing center for COVID
a0_77|NA|drive-thru testing centers for COVID
a0_77|NA|drive-thru testing for COVID
a0_77|NA|drive-thru testing location for COVID
a0_77|NA|drive-thru testing locations for COVID
a0_77|NA|drive-thru testing site for COVID
a0_77|NA|drive-thru testing sites for COVID
a0_77|NA|drive-thru tests for COVID
a0_77|NA|location for a COVID test
a0_77|NA|location for a drive-thru COVID test
a0_77|NA|location for COVID test
a0_77|NA|location for COVID testing
a0_77|NA|location for COVID tests
a0_77|NA|location for drive-thru COVID test
a0_77|NA|location for drive-thru COVID testing
a0_77|NA|location for drive-thru COVID tests
a0_77|NA|locations for a COVID test
a0_77|NA|locations for a drive-thru COVID test
a0_77|NA|locations for COVID test
a0_77|NA|locations for COVID testing
a0_77|NA|locations for COVID tests
a0_77|NA|locations for drive-thru COVID test
a0_77|NA|locations for drive-thru COVID testing
a0_77|NA|locations for drive-thru COVID tests
a0_77|NA|site for a COVID test
a0_77|NA|site for a drive-thru COVID test
a0_77|NA|site for COVID test
a0_77|NA|site for COVID testing
a0_77|NA|site for COVID tests
a0_77|NA|site for drive-thru COVID test
a0_77|NA|site for drive-thru COVID testing
a0_77|NA|site for drive-thru COVID tests
a0_77|NA|sites for a COVID test
a0_77|NA|sites for a drive-thru COVID test
a0_77|NA|sites for COVID test
a0_77|NA|sites for COVID testing
a0_77|NA|sites for COVID tests
a0_77|NA|sites for drive-thru COVID test
a0_77|NA|sites for drive-thru COVID testing
a0_77|NA|sites for drive-thru COVID tests
a0_77|NA|test center for COVID
a0_77|NA|test centers for COVID
a0_77|NA|test for COVID
a0_77|NA|test location for COVID
a0_77|NA|test locations for COVID
a0_77|NA|test site for COVID
a0_77|NA|test sites for COVID
a0_77|NA|tested for COVID
a0_77|NA|testing center for COVID
a0_77|NA|testing centers for COVID
a0_77|NA|testing for COVID
a0_77|NA|testing location for COVID
a0_77|NA|testing locations for COVID
a0_77|NA|testing site for COVID
a0_77|NA|testing sites for COVID
a0_77|NA|tests for COVID
a0_77|NA|center for a drive-through COVID test
a0_77|NA|center for drive-through COVID test
a0_77|NA|center for drive-through COVID testing
a0_77|NA|center for drive-through COVID tests
a0_77|NA|centers for a drive-through COVID test
a0_77|NA|centers for drive-through COVID test
a0_77|NA|centers for drive-through COVID testing
a0_77|NA|centers for drive-through COVID tests
a0_77|NA|COVID drive-through
a0_77|NA|COVID drive-through center
a0_77|NA|COVID drive-through centers
a0_77|NA|COVID drive-through location
a0_77|NA|COVID drive-through locations
a0_77|NA|COVID drive-through site
a0_77|NA|COVID drive-through sites
a0_77|NA|COVID drive-through test
a0_77|NA|COVID drive-through test center
a0_77|NA|COVID drive-through test centers
a0_77|NA|COVID drive-through test location
a0_77|NA|COVID drive-through test locations
a0_77|NA|COVID drive-through test site
a0_77|NA|COVID drive-through test sites
a0_77|NA|COVID drive-through testing
a0_77|NA|COVID drive-through testing center
a0_77|NA|COVID drive-through testing centers
a0_77|NA|COVID drive-through testing location
a0_77|NA|COVID drive-through testing locations
a0_77|NA|COVID drive-through testing site
a0_77|NA|COVID drive-through testing sites
a0_77|NA|COVID drive-through tests
a0_77|NA|drive-through center for a COVID test
a0_77|NA|drive-through center for COVID test
a0_77|NA|drive-through center for COVID testing
a0_77|NA|drive-through center for COVID tests
a0_77|NA|drive-through centers for a COVID test
a0_77|NA|drive-through centers for COVID test
a0_77|NA|drive-through centers for COVID testing
a0_77|NA|drive-through centers for COVID tests
a0_77|NA|drive-through location for a COVID test
a0_77|NA|drive-through location for COVID test
a0_77|NA|drive-through location for COVID testing
a0_77|NA|drive-through location for COVID tests
a0_77|NA|drive-through locations for a COVID test
a0_77|NA|drive-through locations for COVID test
a0_77|NA|drive-through locations for COVID testing
a0_77|NA|drive-through locations for COVID tests
a0_77|NA|drive-through site for a COVID test
a0_77|NA|drive-through site for COVID test
a0_77|NA|drive-through site for COVID testing
a0_77|NA|drive-through site for COVID tests
a0_77|NA|drive-through sites for a COVID test
a0_77|NA|drive-through sites for COVID test
a0_77|NA|drive-through sites for COVID testing
a0_77|NA|drive-through sites for COVID tests
a0_77|NA|drive-through test center for COVID
a0_77|NA|drive-through test centers for COVID
a0_77|NA|drive-through test for COVID
a0_77|NA|drive-through test location for COVID
a0_77|NA|drive-through test locations for COVID
a0_77|NA|drive-through test site for COVID
a0_77|NA|drive-through test sites for COVID
a0_77|NA|drive-through tested for COVID
a0_77|NA|drive-through testing center for COVID
a0_77|NA|drive-through testing centers for COVID
a0_77|NA|drive-through testing for COVID
a0_77|NA|drive-through testing location for COVID
a0_77|NA|drive-through testing locations for COVID
a0_77|NA|drive-through testing site for COVID
a0_77|NA|drive-through testing sites for COVID
a0_77|NA|drive-through tests for COVID
a0_77|NA|location for a drive-through COVID test
a0_77|NA|location for drive-through COVID test
a0_77|NA|location for drive-through COVID testing
a0_77|NA|location for drive-through COVID tests
a0_77|NA|locations for a drive-through COVID test
a0_77|NA|locations for drive-through COVID test
a0_77|NA|locations for drive-through COVID testing
a0_77|NA|locations for drive-through COVID tests
a0_77|NA|site for a drive-through COVID test
a0_77|NA|site for drive-through COVID test
a0_77|NA|site for drive-through COVID testing
a0_77|NA|site for drive-through COVID tests
a0_77|NA|sites for a drive-through COVID test
a0_77|NA|sites for drive-through COVID test
a0_77|NA|sites for drive-through COVID testing
a0_77|NA|sites for drive-through COVID tests
a0_77|NA|center for a drive-by COVID test
a0_77|NA|center for drive-by COVID test
a0_77|NA|center for drive-by COVID testing
a0_77|NA|center for drive-by COVID tests
a0_77|NA|centers for a drive-by COVID test
a0_77|NA|centers for drive-by COVID test
a0_77|NA|centers for drive-by COVID testing
a0_77|NA|centers for drive-by COVID tests
a0_77|NA|COVID drive-by
a0_77|NA|COVID drive-by center
a0_77|NA|COVID drive-by centers
a0_77|NA|COVID drive-by location
a0_77|NA|COVID drive-by locations
a0_77|NA|COVID drive-by site
a0_77|NA|COVID drive-by sites
a0_77|NA|COVID drive-by test
a0_77|NA|COVID drive-by test center
a0_77|NA|COVID drive-by test centers
a0_77|NA|COVID drive-by test location
a0_77|NA|COVID drive-by test locations
a0_77|NA|COVID drive-by test site
a0_77|NA|COVID drive-by test sites
a0_77|NA|COVID drive-by testing
a0_77|NA|COVID drive-by testing center
a0_77|NA|COVID drive-by testing centers
a0_77|NA|COVID drive-by testing location
a0_77|NA|COVID drive-by testing locations
a0_77|NA|COVID drive-by testing site
a0_77|NA|COVID drive-by testing sites
a0_77|NA|COVID drive-by tests
a0_77|NA|drive-by center for a COVID test
a0_77|NA|drive-by center for COVID test
a0_77|NA|drive-by center for COVID testing
a0_77|NA|drive-by center for COVID tests
a0_77|NA|drive-by centers for a COVID test
a0_77|NA|drive-by centers for COVID test
a0_77|NA|drive-by centers for COVID testing
a0_77|NA|drive-by centers for COVID tests
a0_77|NA|drive-by location for a COVID test
a0_77|NA|drive-by location for COVID test
a0_77|NA|drive-by location for COVID testing
a0_77|NA|drive-by location for COVID tests
a0_77|NA|drive-by locations for a COVID test
a0_77|NA|drive-by locations for COVID test
a0_77|NA|drive-by locations for COVID testing
a0_77|NA|drive-by locations for COVID tests
a0_77|NA|drive-by site for a COVID test
a0_77|NA|drive-by site for COVID test
a0_77|NA|drive-by site for COVID testing
a0_77|NA|drive-by site for COVID tests
a0_77|NA|drive-by sites for a COVID test
a0_77|NA|drive-by sites for COVID test
a0_77|NA|drive-by sites for COVID testing
a0_77|NA|drive-by sites for COVID tests
a0_77|NA|drive-by test center for COVID
a0_77|NA|drive-by test centers for COVID
a0_77|NA|drive-by test for COVID
a0_77|NA|drive-by test location for COVID
a0_77|NA|drive-by test locations for COVID
a0_77|NA|drive-by test site for COVID
a0_77|NA|drive-by test sites for COVID
a0_77|NA|drive-by tested for COVID
a0_77|NA|drive-by testing center for COVID
a0_77|NA|drive-by testing centers for COVID
a0_77|NA|drive-by testing for COVID
a0_77|NA|drive-by testing location for COVID
a0_77|NA|drive-by testing locations for COVID
a0_77|NA|drive-by testing site for COVID
a0_77|NA|drive-by testing sites for COVID
a0_77|NA|drive-by tests for COVID
a0_77|NA|location for a drive-by COVID test
a0_77|NA|location for drive-by COVID test
a0_77|NA|location for drive-by COVID testing
a0_77|NA|location for drive-by COVID tests
a0_77|NA|locations for a drive-by COVID test
a0_77|NA|locations for drive-by COVID test
a0_77|NA|locations for drive-by COVID testing
a0_77|NA|locations for drive-by COVID tests
a0_77|NA|site for a drive-by COVID test
a0_77|NA|site for drive-by COVID test
a0_77|NA|site for drive-by COVID testing
a0_77|NA|site for drive-by COVID tests
a0_77|NA|sites for a drive-by COVID test
a0_77|NA|sites for drive-by COVID test
a0_77|NA|sites for drive-by COVID testing
a0_77|NA|sites for drive-by COVID tests
a0_78|NA|COVID-19 testing at home
a0_78|NA|COVID-19 tested at home
a0_78|NA|COVID-19 tests at home
a0_78|NA|COVID-19 test at home
a0_78|NA|at-home COVID-19 testing
a0_78|NA|at-home COVID-19 tested
a0_78|NA|at-home COVID-19 tests
a0_78|NA|at-home COVID-19 test
a0_78|NA|COVID19 testing at home
a0_78|NA|COVID19 tested at home
a0_78|NA|COVID19 tests at home
a0_78|NA|COVID19 test at home
a0_78|NA|at-home COVID19 testing
a0_78|NA|at-home COVID19 tested
a0_78|NA|at-home COVID19 tests
a0_78|NA|at-home COVID19 test
a0_78|NA|COVID testing at home
a0_78|NA|COVID tested at home
a0_78|NA|COVID tests at home
a0_78|NA|COVID test at home
a0_78|NA|at-home COVID testing
a0_78|NA|at-home COVID tested
a0_78|NA|at-home COVID tests
a0_78|NA|at-home COVID test
a0_78|NA|coronavirus testing at home
a0_78|NA|coronavirus tested at home
a0_78|NA|coronavirus tests at home
a0_78|NA|coronavirus test at home
a0_78|NA|at-home coronavirus testing
a0_78|NA|at-home coronavirus tested
a0_78|NA|at-home coronavirus tests
a0_78|NA|at-home coronavirus test
a0_78|NA|COVID-19 testing in home
a0_78|NA|COVID-19 tested in home
a0_78|NA|COVID-19 tests in home
a0_78|NA|COVID-19 test in home
a0_78|NA|in-home COVID-19 testing
a0_78|NA|in-home COVID-19 tested
a0_78|NA|in-home COVID-19 tests
a0_78|NA|in-home COVID-19 test
a0_78|NA|COVID19 testing in home
a0_78|NA|COVID19 tested in home
a0_78|NA|COVID19 tests in home
a0_78|NA|COVID19 test in home
a0_78|NA|in-home COVID19 testing
a0_78|NA|in-home COVID19 tested
a0_78|NA|in-home COVID19 tests
a0_78|NA|in-home COVID19 test
a0_78|NA|COVID testing in home
a0_78|NA|COVID tested in home
a0_78|NA|COVID tests in home
a0_78|NA|COVID test in home
a0_78|NA|in-home COVID testing
a0_78|NA|in-home COVID tested
a0_78|NA|in-home COVID tests
a0_78|NA|in-home COVID test
a0_78|NA|coronavirus testing in home
a0_78|NA|coronavirus tested in home
a0_78|NA|coronavirus tests in home
a0_78|NA|coronavirus test in home
a0_78|NA|in-home coronavirus testing
a0_78|NA|in-home coronavirus tested
a0_78|NA|in-home coronavirus tests
a0_78|NA|in-home coronavirus test
a0_79|NA|COVID-19 signs and symptoms
a0_79|NA|COVID-19 symptoms
a0_79|NA|sign of COVID-19
a0_80|NA|rule-out COVID-19
a0_80|NA|rule-out COVID19
a0_80|NA|rule-out COVID
a0_80|NA|rule-out the novel coronavirus
a0_80|NA|rule-out novel coronavirus
a0_80|NA|r/o COVID-19
a0_80|NA|r/o COVID19
a0_80|NA|r/o COVID
a0_80|NA|r/o the novel coronavirus
a0_80|NA|r/o novel coronavirus
a0_81|NA|public health emergency
a0_81|NA|public health emergencies
a0_81|NA|public health crisis
a0_81|NA|public health crises
a0_81|NA|health emergency
a0_81|NA|health emergencies
a0_81|NA|health crisis
a0_81|NA|health crises
a0_82|NA|COVID-19 test
a0_82|NA|COVID-19 testing
a0_82|NA|COVID-19 tests
a0_82|NA|testing for COVID-19
a0_82|NA|tested for COVID-19
a0_82|NA|tests for COVID-19
a0_82|NA|test for COVID-19
a0_82|NA|testing COVID-19
a0_82|NA|tested COVID-19
a0_82|NA|tests COVID-19
a0_82|NA|test COVID-19
a0_82|NA|COVID19 test
a0_82|NA|COVID19 tested
a0_82|NA|COVID19 testing
a0_82|NA|COVID19 tests
a0_82|NA|testing for COVID19
a0_82|NA|tested for COVID19
a0_82|NA|tests for COVID19
a0_82|NA|test for COVID19
a0_82|NA|testing COVID19
a0_82|NA|tested COVID19
a0_82|NA|tests COVID19
a0_82|NA|test COVID19
a0_82|NA|COVID test
a0_82|NA|COVID testing
a0_82|NA|COVID tests
a0_82|NA|testing for COVID
a0_82|NA|tested for COVID
a0_82|NA|tests for COVID
a0_82|NA|test for COVID
a0_82|NA|testing COVID
a0_82|NA|tested COVID
a0_82|NA|tests COVID
a0_82|NA|test COVID
a0_82|NA|coronavirus test
a0_82|NA|coronavirus testing
a0_82|NA|coronavirus tests
a0_82|NA|testing for coronavirus
a0_82|NA|tested for coronavirus
a0_82|NA|tests for coronavirus
a0_82|NA|test for coronavirus
a0_82|NA|testing coronavirus
a0_82|NA|tested coronavirus
a0_82|NA|test coronavirus
a0_82|NA|tests coronavirus
a0_82|NA|novel coronavirus test
a0_82|NA|novel coronavirus testing
a0_82|NA|novel coronavirus tests
a0_82|NA|testing for novel coronavirus
a0_82|NA|tested for novel coronavirus
a0_82|NA|tests for novel coronavirus
a0_82|NA|test for novel coronavirus
a0_82|NA|testing novel coronavirus
a0_82|NA|tested novel coronavirus
a0_82|NA|tests novel coronavirus
a0_82|NA|test novel coronavirus
a0_82|NA|new coronavirus test
a0_82|NA|new coronavirus testing
a0_82|NA|new coronavirus tests
a0_82|NA|testing for new coronavirus
a0_82|NA|tested for new coronavirus
a0_82|NA|tests for new coronavirus
a0_82|NA|test for new coronavirus
a0_82|NA|testing new coronavirus
a0_82|NA|tested new coronavirus
a0_82|NA|tests new coronavirus
a0_82|NA|test new coronavirus
a0_82|NA|tested for the coronavirus
a0_82|NA|tested for the new coronavirus
a0_82|NA|tested for the novel coronavirus
a0_82|NA|testing for the coronavirus
a0_82|NA|testing for the new coronavirus
a0_82|NA|testing for the novel coronavirus
a0_82|NA|tests for the coronavirus
a0_82|NA|test for the coronavirus
a0_82|NA|tests for the new coronavirus
a0_82|NA|test for the new coronavirus
a0_82|NA|tests for the novel coronavirus
a0_82|NA|test for the novel coronavirus
a0_83|NA|hydroxychloroquine sulfate
a0_83|NA|hydroxychloroquine
a0_83|NA|hydroxy-chloroquine sulfate
a0_83|NA|hydroxy-chloroquine
a0_83|NA|HCQ
a0_84|NA|full face mask
a0_84|NA|FFM
a0_84|NA|face mask
a0_84|NA|full face masks
a0_84|NA|FFMs
a0_84|NA|face masks
a0_85|NA|PUI
a0_85|NA|person under investigation
a0_86|NA|COVID-19 signs and symptoms
a0_86|NA|COVID-19 signs
a0_86|NA|sign of COVID-19
BMV_1|C0220781|Anabolism
BMV_2|NA|antibody response
BMV_3|NA|antiviral
BMV_3|NA|antivirals
BMV_4|NA|antiviral activity
BMV_4|NA|antiviral activities
BMV_5|C0003451|Antiviral Agents
BMV_6|C0162638|Apoptosis
BMV_7|C0004391|Autophagy
BMV_8|NA|B-cell assays
BMV_9|NA|B-cell epitopes
BMV_10|C0004793|Base Sequence
BMV_11|C0005507|Biological Assay
BMV_12|C0005528|Biological Transport
BMV_13|NA|bronchoalveolar lavage fluid
BMV_13|NA|BALF
BMV_14|C0007584|Cell Count
BMV_15|C0007587|Cell Death
BMV_16|C0007589|Cell Differentiation process
BMV_17|C0007609|Cell Nucleolus
BMV_18|NA|chest radiography
BMV_19|NA|clinical characteristic
BMV_19|NA|clinical characteristics
BMV_20|NA|clinical data
BMV_20|NA|clinical datas
BMV_21|NA|clinical experimental vaccine research
BMV_22|NA|clinical importance
BMV_23|NA|clinical sign
BMV_23|NA|clinical signs
BMV_24|C0008972|Clinical Study
BMV_25|NA|confirmed cas
BMV_25|NA|confirmed cases
BMV_26|NA|conformational masking
BMV_27|NA|cross-neutralization
BMV_28|NA|cross-neutralizing antibody
BMV_28|NA|cross-neutralizing antibodies
BMV_29|NA|Cryo-EM structure
BMV_30|C1511760|Deletion Mutation
BMV_31|C0011900|diagnosis
BMV_31|C0011900|diagnoses
BMV_32|C0242781|disease transmission
BMV_33|C0598312|DNA Replication
BMV_34|C0162326|DNA Sequence
BMV_35|C0013220|Drug Tolerance
BMV_36|C2745965|Emergencies
BMV_36|C2745965|emergency
BMV_37|C0014441|Enzyme-Linked Immunosorbent Assay
BMV_37|C0014441|elisa
BMV_38|C0014507|Epidemiology
BMV_39|NA|epitope
BMV_39|NA|epitopes
BMV_40|NA|fecal sample
BMV_40|NA|fecal samples
BMV_41|C0017262|Gene Expression
BMV_42|C0017296|Gene therapy
BMV_43|C0017337|Genes
BMV_43|C0017337|gene
BMV_44|C0042333|Genetic Diversity
BMV_45|C0034865|Genetic Recombination
BMV_46|C0036576|Genetic Selection
BMV_47|C0040649|Genetic Transcription
BMV_48|C0017428|Genome
BMV_49|C1456573|Global Health
BMV_50|NA|global pandemic
BMV_51|NA|glycan shielding
BMV_52|NA|glycoprotein
BMV_52|NA|glycoproteins
BMV_53|C0677043|histopathology
BMV_54|NA|homotrimer
BMV_54|NA|homotrimers
BMV_55|NA|host cell
BMV_55|NA|host cells
BMV_56|C0020517|Hypersensitivity
BMV_57|NA|immune cell
BMV_57|NA|immune cells
BMV_58|NA|immune response
BMV_58|NA|immune responses
BMV_59|C0020963|Immune Tolerance
BMV_60|C0020971|Immunization
BMV_61|NA|immunoblotting
BMV_62|NA|immunofluorescence test
BMV_63|NA|immunogenicity
BMV_64|NA|immunolobulin g
BMV_64|NA|igg
BMV_65|NA|incubation period
BMV_65|NA|incubation periods
BMV_66|NA|induction
BMV_67|NA|infectivity
BMV_68|NA|inhibition
BMV_68|NA|inhibitions
BMV_69|NA|interaction
BMV_69|NA|interactions
BMV_70|C0220862|isolation
BMV_71|NA|low-input metagenomic next-generation sequencing
BMV_71|NA|mNGS
BMV_72|NA|lungs
BMV_73|C0024432|"Macrophage | macrophages"
BMV_74|NA|Major histocompatibility complex binding assays
BMV_75|C2936622|Massively-Parallel Sequencing
BMV_76|C0199470|Mechanical Ventilation
BMV_77|C0025246|Membrane Fusion
BMV_78|NA|MHC binding assays
BMV_79|NA|microbiol
BMV_80|NA|molecular mechanisms
BMV_81|C0220880|morbidity
BMV_82|C0026882|Mutation
BMV_82|C0026882|mutations
BMV_83|NA|nasopharyngeal swabs
BMV_84|NA|next-generation sequencing
BMV_84|NA|ngs
BMV_85|NA|nucleolus
BMV_86|C0206415|Oligonucleotide Primers
BMV_87|NA|orf
BMV_88|NA|overexpression
BMV_89|NA|pathogen
BMV_89|NA|pathogens
BMV_90|NA|pathogenicity
BMV_91|C1136169|Pathogenicity
BMV_92|C0030657|pathogenicity
BMV_93|NA|pathway
BMV_93|NA|pathways
BMV_94|C0013227|Pharmaceutical Preparations
BMV_95|C0013216|Pharmacotherapy
BMV_96|C0031715|Phosphorylation
BMV_97|NA|primer
BMV_97|NA|primers
BMV_98|C0184661|Procedures
BMV_99|C0033613|Protective Agents
BMV_100|C0597295|Protein Biosynthesis
BMV_101|NA|protein expression
BMV_102|C0034019|Public Health
BMV_103|C0243114|purification
BMV_104|NA|recombination
BMV_105|NA|replication
BMV_106|C0035168|Research
BMV_107|C0242481|Research Activities
BMV_108|C0035171|Research Design
BMV_109|NA|respiratory infection
BMV_109|NA|respiratory infections
BMV_110|C0599161|Reverse Transcriptase Polymerase Chain Reaction
BMV_110|C0599161|rt-pcr
BMV_111|NA|RNA analysis
BMV_112|C1136031|RNA Interference
BMV_112|C1136031|rnai
BMV_113|C1522002|RNA Recognition Motif
BMV_114|C0162327|RNA Sequence
BMV_115|NA|RNA virus
BMV_116|NA|rnvirus
BMV_116|NA|rnviruses
BMV_117|NA|sequence
BMV_117|NA|sequences
BMV_118|C0162801|Sequence Analysis
BMV_119|NA|serum
BMV_119|NA|sera
BMV_120|C0752046|Single Nucleotide Polymorphism
BMV_120|C0752046|snp
BMV_120|C0752046|snps
BMV_120|C0752046|single nucleotide polymorphisms
BMV_121|C0220921|survival
BMV_122|C0683368|symptoms
BMV_123|NA|T-cell assays
BMV_124|NA|T-cell epitopes
BMV_125|C0087111|Therapeutics
BMV_126|C0039798|therapy
BMV_127|C3665494|Thoracic Radiography
BMV_128|NA|transcription
BMV_129|NA|transfection
BMV_129|NA|transfections
BMV_130|NA|transmissibility
BMV_131|C0042196|Vaccination
BMV_132|NA|vaccine design
BMV_133|NA|viral entry
BMV_134|C0035736|Viral RNA
BMV_135|C0042765|Virulence
BMV_136|C0220936|virulence
BMV_137|C1537068|Virus Internalization
BMV_138|C0042774|Virus Replication
BMV_138|C0042774|virus replications
BMV_138|C0042774|viral replication
BMV_138|C0042774|viral replications
BMV_139|NA|Western-Blot
BMV_139|NA|western-blotting
BMV_139|NA|WB
BMV_139|NA|Western-Blot
BMV_139|NA|western-blotting
BMV_139|NA|WB
CL_1|NA|Caco-2
CL_2|NA|Calu-3
CL_3|NA|Calu-3 2B4
CL_4|NA|HEK293T
CL_4|NA|293T 
CL_5|NA|Huh-7
CL_6|NA|Vero
CL_7|NA|VeroE6
CL_7|NA|Vero C1008
CL_8|NA|VeroE6/TMPRSS2
CL_9|NA|CHO-K1
CL_10|NA|K-562
CL_11|NA|PER.C6
CL_12|NA|47D11
CL_13|NA|F26G1
CL_14|NA|F26G6
CL_15|NA|F26G8
CL_16|NA|F26G18
CL_17|NA|F26G19
CL_18|NA|N-176-15
CL_19|NA|S-9-11
CL_20|NA|rSN-18
CL_21|NA|rSN-21-2
CL_22|NA|rSN-29
CL_23|NA|rSN-122
CL_24|NA|rSN-150
DG_1|NA|Acetylcysteine
DG_1|NA|"Acetadote | Cetylev | Mucomyst | Parvolex"
DG_2|NA|Adalimumab
DG_3|NA|Amprenavir
DG_3|NA|(3S)-Tetrahydro-3-furanyl ((1S,2R)-3-(((4-aminophenyl)sulfonyl)(2-methylpropyl)amino)-2-hydroxy-1-(phenylmethyl)propyl)carbamate
DG_4|NA|Angiotensin II
DG_28|NA|Artenimol
DG_28|NA|Dihydroartemisinin
DG_7|NA|ASC09
DG_5|NA|Atazanavir
DG_5|NA|"Reyataz | Atavir | ATZ"
DG_6|NA|Atovaquone
DG_6|NA|2-(trans-4-(p-Chlorophenyl)cyclohexyl)-3-hydroxy-1,4-naphthoquinone
DG_8|NA|Aviptadil
DG_8|NA|RLF-100
DG_9|NA|Azithromycin
DG_9|NA|AzaSite
DG_10|NA|Azvudine
DG_10|NA|RO-0622
DG_11|NA|Baloxavir marboxil
DG_11|NA|Xofluza
DG_12|NA|Baricitinib
DG_12|NA|Olumiant
DG_13|NA|Bepotastine
DG_13|NA|Bepreve
DG_14|NA|Bismuth potassium citrate
DG_14|NA|Pylera
DG_15|NA|Bromhexine hydrochloride
DG_15|NA|Bisolvon
DG_16|NA|Camrelizumab
DG_17|NA|Carriomycin
DG_18|NA|CD24Fc
DG_19|NA|Cefditoren
DG_19|NA|Spectracef
DG_20|NA|Cefixime
DG_20|NA|Suprax
DG_21|C0008269|Chloroquine
DG_21|C0008269|Nivaquine
DG_21|C0008269|N4-(7-chloro-4-quinolinyl)-N1,N1-diethyl-1,4-pentanediamine
DG_22|NA|Clarithromycin
DG_22|NA|"6-O-methyl erythromycin | Biaxin"
DG_23|NA|Cobicistat
DG_23|NA|Tybost
DG_24|NA|Danoprevir
DG_24|NA|Ganovo
DG_25|NA|Darunavir
DG_25|NA|Prezista
DG_26|NA|Daunorubicin
DG_26|NA|Cerubidine
DG_27|NA|Diammonium glycyrrhizinate
DG_29|NA|Dipyridamole
DG_29|NA|"Agilease | Cardoxin | Cleridium"
DG_29|NA|Curantyl
DG_29|NA|Persantin
DG_30|NA|Ebastine
DG_31|NA|Eculizumab
DG_31|NA|Soliris
DG_32|NA|Erythromycin
DG_32|NA|Abomacetin
DG_32|NA|Ilosone
DG_33|NA|Favipiravir
DG_33|NA|"Avigan | T-705"
DG_34|NA|Fingolimod
DG_34|NA|"Gilenya | Gilenia"
DG_35|NA|Fosamprenavir
DG_35|NA|FOS-APV
DG_36|NA|Galidesivir
DG_36|NA|Immucillin A
DG_37|NA|Hydrogen peroxide
DG_37|NA|Eskata
DG_38|NA|Hydroxychloroquine
DG_38|NA|Oxichloroquine
DG_38|NA|"Oxichlorochine | Plaquenil | Dolquine | HCQS | Quensyl"
DG_38|NA|Polirreumin
DG_78|NA|ibuprofen
DG_39|NA|Indinavir
DG_39|NA|Crixivan
DG_40|NA|Inhaled gases
DG_41|NA|Interferon alfacon-1
DG_41|NA|"IFN Alfacon-1 | IFN-Con1 | Interferon alfacon-1 | Infergen"
DG_42|NA|Ivermectin
DG_42|NA|"Stromectol | Ascapil"
DG_42|NA|"Detebencil | Ermetin | Gotax"
DG_42|NA|Imectin
DG_42|NA|Ivectin
DG_42|NA|Ivera
DG_42|NA|Ivergot
DG_42|NA|Ivermec
DG_42|NA|Ivexterm
DG_42|NA|Ivori
DG_42|NA|Kaonol
DG_42|NA|Kilox
DG_42|NA|Maikeding
DG_42|NA|Quanox
DG_42|NA|Revectina
DG_42|NA|Scabo
DG_42|NA|Scavista
DG_42|NA|Securo
DG_42|NA|Vermectin
DG_43|NA|Jakotinib hydrochloride
DG_44|NA|Leflunomide
DG_44|NA|Arava
DG_45|NA|Lopinavir
DG_45|NA|Kaletra
DG_79|NA|marijuana
DG_46|NA|Mepolizumab
DG_46|NA|Nucala
DG_47|NA|Metamizole
DG_47|NA|Algocalmin
DG_47|NA|Algozone
DG_47|NA|Analgin
DG_47|NA|Dimethone
DG_47|NA|Dipirona
DG_47|NA|Neo-Melubrina
DG_47|NA|Novalgin
DG_47|NA|Optalgin
DG_47|NA|Protemp
DG_47|NA|Pyralgin
DG_48|NA|Methylprednisolone
DG_48|NA|"Depo-Medrol | Hybrisil | Medrol | Medroloan"
DG_49|NA|Mitoxantrone
DG_49|NA|Novantrone
DG_50|NA|Moexipril
DG_50|NA|Univasc
DG_51|NA|MSCs
DG_52|NA|Nelfinavir
DG_52|NA|Viracept
DG_53|NA|NestCell®
DG_54|NA|PD-1 mAb
DG_54|NA|PD1
DG_54|NA|PD-1
DG_54|NA|PD1 mAb
DG_80|NA|penicillin
DG_55|NA|Pirfenidone
DG_55|NA|Esbriet
DG_56|NA|Polyinosinic-polycytidylic acid
DG_57|NA|PUL-042 Inhalation Solution
DG_58|NA|Remdesivir
DG_58|NA|GS-5734
DG_59|NA|rhG-CSF
DG_60|NA|Ribavirin
DG_61|NA|Ritonavir
DG_61|NA|Norvir
DG_62|NA|Rosuvastatin
DG_62|NA|Crestor
DG_63|NA|Ruxolitinib
DG_63|NA|"Jakafi | Jakavi"
DG_64|NA|Saquinavir
DG_64|NA|Invirase
DG_65|NA|Sarilumab
DG_66|NA|Sildenafil
DG_67|NA|Sofosbuvir
DG_67|NA|Sovaldi
DG_68|NA|Suramin sodium
DG_69|NA|Thalidomide
DG_69|NA|Thalomid
DG_70|NA|Thymosin
DG_71|NA|Tipranavir
DG_71|NA|Aptivus
DG_72|NA|Tocilizumab
DG_72|NA|"Actemra | Atlizumab"
DG_73|NA|Tranilast
DG_74|NA|Triazavirin
DG_75|NA|UC-MSCs
DG_76|NA|Umifenovir
DG_76|NA|"Arbidol | Arbidole"
DG_77|NA|Vitamin C
CE_1|NA|“crown-like” appearance
CE_2|C0206132|age of onset
CE_3|C1524024|analysis
CE_4|NA|antiserum
CE_4|NA|antisera
CE_5|C0243073|assay
CE_6|NA|astrovirus
CE_6|NA|astroviruses
CE_7|NA|asymptomatic
CE_7|NA|asymptomatical
CE_8|NA|cluster
CE_8|NA|clusters
CE_9|NA|contact tracing
CE_10|NA|containment
CE_11|NA|contamination
CE_11|NA|contaminations
CE_12|C0243148|control
CE_13|NA|control measure
CE_13|NA|control measures
CE_14|NA|coronavirus
CE_14|NA|coronaviruses
CE_15|NA|crucial role
CE_15|NA|crucial roles
CE_16|NA|cumulative number
CE_16|NA|cumulative numbers
CE_17|NA|current study
CE_17|NA|current studies
CE_18|C0993637|Database
CE_19|C0011065|Death
CE_20|C0011750|Developing Countries
CE_20|C0011750|developing country
CE_21|NA|diabete
CE_22|NA|diagnosis
CE_23|C1704711|distribution
CE_24|NA|emergency
CE_24|NA|emergencies
CE_25|NA|epicenter
CE_26|C0220823|epidemics
CE_26|C0220823|epidemic
CE_27|NA|epidemiological investigation
CE_27|NA|epidemiological investigations
CE_28|NA|epidemiology
CE_29|NA|expression level
CE_29|NA|expression levels
CE_30|C2607943|findings
CE_31|C0815319|Geographic Information Systems
CE_32|C0017446|Geographic Locations
CE_33|C0220844|growth
CE_34|C0282423|Guideline
CE_35|C0162791|Guidelines
CE_36|C0220845|guiding characteristics
CE_37|NA|health emergency
CE_37|NA|health emergencies
CE_38|C0018724|Health Personnel
CE_39|NA|healthcare workers
CE_39|NA|health care workers
CE_40|NA|hospitalisation
CE_41|NA|host
CE_42|NA|Huanan market
CE_42|NA|Huanan markets
CE_43|NA|human health
CE_44|NA|human-to-human transmission
CE_45|NA|immune response
CE_45|NA|immune responses
CE_46|NA|immunity
CE_47|NA|imported case
CE_47|NA|imported cases
CE_48|C0220856|incidence
CE_49|NA|incubation period
CE_49|NA|incubation periods
CE_50|NA|infected animal
CE_50|NA|infected animals
CE_51|NA|intermediate host
CE_51|NA|intermediate hosts
CE_52|NA|international concern
CE_53|NA|large number
CE_53|NA|large numbers
CE_54|NA|lethality
CE_55|C0876936|Mathematical Model
CE_55|C0876936|mathematical models
CE_56|C0025106|Medical Staff
CE_57|C0025266|Men
CE_58|C0026565|Mortality
CE_59|C0026566|mortality
CE_60|NA|nasopharyngeal sample
CE_60|NA|nasopharyngeal samples
CE_61|NA|oropharyngeal sample
CE_61|NA|oropharyngeal samples
CE_62|NA|oxygen
CE_63|C1615608|Pandemics
CE_63|C1615608|pandemic
CE_64|NA|patient
CE_64|NA|patients
CE_65|NA|permission
CE_65|NA|permissions
CE_66|C0031166|Permissiveness
CE_67|NA|person-to-person transmission
CE_68|C0031843|physiology
CE_69|C0032659|Population
CE_70|C1257890|Population Group
CE_71|NA|positive rate
CE_72|NA|preparedness
CE_73|C0033105|Prevalence
CE_74|C0220900|prevalence
CE_75|C2700409|prevention
CE_76|NA|public health emergency
CE_77|NA|public health emergency of international concern
CE_78|NA|publicly funded repository
CE_78|NA|publicly funded repositories
CE_79|NA|quarantine
CE_80|C0035173|Research Personnel
CE_81|C0035648|Risk Factors
CE_81|C0035648|risk factor
CE_82|C0035691|RNA Viruses
CE_82|C0035691|rna virus
CE_83|NA|rnvirus
CE_83|NA|rnviruses
CE_84|NA|school closures
CE_85|C0036667|Sensitivity
CE_86|NA|serum
CE_86|NA|sera
CE_87|C1522384|Sex
CE_88|NA|shortness of breath
CE_89|C0037412|Social Distance
CE_89|C0037412|social distancing
CE_90|C0037791|Specificity
CE_91|NA|study design
CE_92|NA|subset
CE_93|NA|supplementary information
CE_94|C0220920|surveillance
CE_95|C0040722|transmission
CE_96|C0040802|Travel
CE_97|NA|treatment
CE_98|NA|trimer
CE_98|NA|trimers
CE_99|NA|urgent need
CE_100|NA|vaccination
CE_100|NA|vaccinations
CE_101|NA|vaccine
CE_101|NA|vaccines
CE_102|NA|vast majority
CE_103|NA|vector-born
CE_104|C0242856|Veterinarian
CE_105|C0521026|viruses
CE_105|C0521026|virus
CE_106|NA|wide range
CE_107|NA|World Health Organization
CE_107|NA|WHO
CE_108|NA|zoonose
CE_109|C1552907|Adenovirus Vaccine
DIS_1|NA|abdominal pain
DIS_2|NA|acetaminophen
DIS_3|NA|acute respiratory distress syndrome
DIS_3|NA|"ARDS | respiratory distress"
DIS_4|NA|afebrile
DIS_5|NA|albuterol
DIS_6|NA|anaphylaxis
DIS_7|NA|anemia
DIS_8|NA|anxiety
DIS_9|NA|asthma
DIS_10|NA|chest pain
DIS_11|NA|chills
DIS_12|C0024117|Chronic Obstructive Airway Disease
DIS_13|NA|Chronic obstructive pulmonary disease
DIS_13|NA|copd
DIS_14|C0275524|Coinfection
DIS_15|C0009450|Communicable Diseases
DIS_16|NA|congestion
DIS_18|C0206750|Coronavirus Infections
DIS_19|C0010200|cough
DIS_19|C0010200|Coughing
DIS_20|NA|depression
DIS_21|NA|diabete
DIS_21|NA|diabetes
DIS_22|NA|diarrhea
DIS_23|NA|diffuse alveolar damage
DIS_24|NA|dry cough
DIS_25|NA|dyspnea
DIS_26|NA|edema
DIS_27|C0872315|Emerging Communicable Diseases
DIS_28|NA|emerging infectious disease
DIS_28|NA|emerging infectious diseases
DIS_29|NA|fatigue
DIS_30|NA|febrile
DIS_31|NA|fever
DIS_32|NA|gastroesophageal reflux disorder
DIS_33|NA|headache
DIS_34|NA|hyperlipidemia
DIS_35|NA|hypertension
DIS_36|NA|infection
DIS_36|NA|infections
DIS_37|NA|infectious disease
DIS_37|NA|infectious diseases
DIS_38|NA|influenza
DIS_39|NA|malaise
DIS_40|NA|mers-cov infection
DIS_41|C3694279|Middle East Respiratory Syndrome
DIS_41|C3694279|MERS
DIS_42|NA|myalgia
DIS_43|NA|nausea
DIS_44|NA|vomiting
DIS_45|NA|nausea and vomiting
DIS_46|NA|Novel Coronavirus Pneumonia
DIS_46|NA|ncp
DIS_48|NA|pain
DIS_50|NA|pneumonia
DIS_51|NA|pruritis
DIS_51|NA|itchy skin
DIS_51|NA|pruritus
DIS_52|NA|rales
DIS_52|NA|crackles
DIS_53|NA|rash
DIS_54|NA|respiratory disease
DIS_54|NA|respiratory diseases
DIS_55|C0035222|Respiratory Distress Syndrome
DIS_56|NA|respiratory infection
DIS_56|NA|respiratory infections
DIS_57|C0035243|Respiratory Tract Infections
DIS_58|NA|rhinorrhea
DIS_59|NA|sepsis
DIS_60|C1175175|Severe Acute Respiratory Syndrome
DIS_60|C1175175|SARS
DIS_61|NA|sore throat
DIS_62|NA|sputum
DIS_63|NA|sulfonamide antibiotic
DIS_63|NA|sulfonamide antibiotics
DIS_64|NA|tachycardia
DIS_65|NA|tachypnea
DIS_66|NA|urticaria
DIS_67|NA|viral illness
DIS_68|NA|viral respiratory infection
DIS_68|NA|viral respiratory infections
DIS_69|C0042769|Virus Diseases
DIS_70|NA|virus infection
DIS_70|NA|virus infections
DIS_70|NA|viral infection
DIS_70|NA|viral infections
DIS_71|NA|weakness
DIS_72|NA|wheezing
SP_1|C2806453|Betacoronavirus
SP_2|C0006801|Camel
SP_2|C0006801|camels
SP_3|C0013127|Camelus dromedarius
SP_3|C0013127|dromedary
SP_3|C0013127|dromaderies
SP_4|C0206419|Coronavirus
SP_4|C0206419|coronaviruses
SP_4|C0206419|cov
SP_4|C0206419|covs
SP_5|NA|COVID-19
SP_5|NA|Severe Acute Respiratory Syndrome Coronavirus 2
SP_5|NA|SARS-CoV-2
SP_5|NA|2019-nCoV
SP_6|C1510418|dog
SP_6|C1510418|canis lupus
SP_7|NA|dromedary camels
SP_7|NA|dromedary camel
SP_8|C4168815|HKU23
SP_8|C4168815|Camel coronavirus HKU23
SP_9|C0086418|Homo sapiens
SP_9|C0086418|Human
SP_10|C0206422|human coronavirus
SP_10|C0206422|hcov
SP_11|C4316910|influenza virus
SP_11|C4316910|influenzvirus
SP_12|C3698360|MERS-CoV
SP_12|C3698360|"Middle East Respiratory Syndrome Coronavirus | MERS Coronavirus"
SP_13|NA|novel coronavirus
SP_14|C0325072|Paguma larvata
SP_14|C0325072|"Palm civet | Paradoxurus hermaphroditus"
SP_14|C0325072|"palm civets | Masked palm civet"
SP_15|C0999626|Manidae
SP_15|C0999626|pangolin
SP_15|C0999626|pangolins
SP_16|C0597404|respiratory viruses
SP_17|C1218105|Rhinolophus macrotis
SP_17|C1218105|"Horseshoe bats | Rhinolophus | Big-eared horseshoe bat"
SP_18|C1175743|SARS-CoV
SP_18|C1175743|"Severe acute respiratory distress syndrome coronavirus | SARS coronavirus"
SP_19|C0008139|Chiroptera
SP_19|C0008139|bat
SP_19|C0008139|bats
SP_20|C1676985|HKU1
SP_20|C1676985|Human coronavirus HKU1
SP_21|C0949881|OC43
SP_21|C0949881|Human coronavirus OC43
PG_1|NA|3cl pro
PG_2|C1422064|ACE2
PG_3|C1452534|Angiontensin-converting enyme human protein
PG_3|C1452534|ACE human protein
PG_4|C1610422|Angiotensin-converting enzyme 2
PG_4|C1610422|"hACE2 | human ACE2 | ACE2 | human Angiotensin-converting enzyme 2 | ACE-related carboxypeptidase | ACEH "
PG_5|C0003018|Angiotensins
PG_6|C0966484|CLEC4M
PG_6|C0966484|C-type lectin domain family 4 member M
PG_7|C1539099|CLEC4M
PG_7|C1539099|CD209L
PG_8|C0079189|Cytokines
PG_8|C0079189|cytokine
PG_9|C1447020|DPP4
PG_9|C1447020|CD26
PG_10|C1414141|DPP4
PG_11|NA|Envelope small membrane protein
PG_11|NA|"E protein | small enveloppe protein | sM protein"
PG_12|NA|interferon
PG_12|NA|ifn
PG_13|C0085295|Interleukin-10
PG_13|C0085295|il-10
PG_14|C1699802|IL10 human protein
PG_15|NA|matrix protein
PG_15|NA|M protein
PG_16|C0003250|Monoclonal Antibodies
PG_17|C0475463|Neutralizing Antibodies
PG_17|C0475463|neutralizing antibody
PG_18|NA|Nucleoprotein
PG_18|NA|"N protein | nucleocapsid protein "
PG_19|C0033382|Proline
PG_20|NA|Protein 3a
PG_20|NA|"Protein U274 | Protein X1"
PG_21|NA|Protein 7a
PG_21|NA|"Accessory protein 7a | Protein U122"
PG_21|NA|Protein X4
PG_22|NA|Replicase polyprotein 1a
PG_23|NA|Replicase polyprotein 1a
PG_23|NA|pp1a
PG_24|NA|Replicase polyprotein 1ab
PG_25|NA|Replicase polyprotein 1ab
PG_25|NA|pp1ab
PG_26|NA|RNA-dependent RNA polymerase
PG_26|NA|rdrp
PG_26|NA|rdr
PG_26|NA|RNA replicase
PG_27|NA|SARS-CoV-2 RBD
PG_28|C3711684|SARS-S
PG_29|NA|Spike glycoprotein
PG_29|NA|S protein
PG_29|NA|"Spike glycoprotein | Peplomer protein | E2"
PG_30|NA|Spike glycoprotein
PG_30|NA|S glycoprotein
PG_31|NA|TMPRSS2
PG_31|NA|PRSS10
PG_32|NA|Transmembrane protease serine 2
PG_32|NA|Serine protease 10
