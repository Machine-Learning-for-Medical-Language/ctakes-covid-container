##  Columns = CUI|TUI|STR|PREF
C0027424|T184|nasal congestion|Congestion or runny nose
C0027424|T184|stuffed-up nose|Congestion or runny nose
C0027424|T184|stuffy nose|Congestion or runny nose
C0027424|T184|congested nose|Congestion or runny nose
C1260880|T184|rhinorrhea|Congestion or runny nose
C1260880|T184|Nasal discharge|Congestion or runny nose
C1260880|T184|discharge from nose|Congestion or runny nose
C1260880|T184|nose dripping|Congestion or runny nose
C1260880|T184|nose running|Congestion or runny nose
C1260880|T184|running nose|Congestion or runny nose
C1260880|T184|runny nose|Congestion or runny nose
C0027424|T184|R09.81|Congestion or runny nose
C0010200|T184|cough|Cough
C0010200|T184|coughing|Cough
C0010200|T184|tussive|Cough
C0010200|T184|posttussive|Cough
C0010200|T184|post-tussive|Cough
C0010200|T184|R05|Cough
C0010200|T184|R05.9|Cough
C0850149|T184|dry cough|Cough
C0850149|T184|dry coughs|Cough
C0850149|T184|coughs dry|Cough
C0850149|T184|unproductive cough|Cough
C0850149|T184|non-productive cough|Cough
C0239134|T033|productive cough|Cough
C0239134|T033|loose cough|Cough
C0239134|T033|moist cough|Cough
C0239134|T033|Producing sputum|Cough
C0239134|T033|Bronchial cough|Cough
C0239134|T033|Chest cough|Cough
C0239134|T033|Chesty cough|Cough
C0011991|T184|diarrhea|Diarrhea
C0011991|T184|R19.7|Diarrhea
C0011991|T184|Watery stool|Diarrhea
C0011991|T184|Watery stools|Diarrhea
C0015672|T184|fatigue|Fatigue
C0015672|T184|fatigues|Fatigue
C0015672|T184|fatigued|Fatigue
C0015672|T184|tiredness|Fatigue
C0015672|T184|lack of energy|Fatigue
C0015672|T184|energy loss|Fatigue
C0015672|T184|weariness|Fatigue
C0015672|T184|R53.83|Fatigue
C0231218|T184|Malaise|Fatigue
C0231218|T184|Generally unwell|Fatigue
C0231218|T184|R53.81|Fatigue
C0085593|T184|Chill|Fever or chills
C0085593|T184|Chills|Fever or chills
C0085593|T184|R68.83|Fever or chills
C0015967|T184|Fever|Fever or chills
C0015967|T184|Fevers|Fever or chills
C0015967|T184|Pyrexia|Fever or chills
C0085594|T184|Fever with chills|Fever or chills
C0085594|T184|Fever and chills|Fever or chills
C0085594|T184|Pyrexia with chills|Fever or chills
C0085594|T184|Fever Chills|Fever or chills
C0085594|T184|R50|Fever or chills
C0085594|T184|R50.0|Fever or chills
C0085594|T184|R50.9|Fever or chills
C0018681|T184|Headache|Headache
C0018681|T184|HA|Headache
C0018681|T184|Cephalgia|Headache
C0018681|T184|Cephalalgia|Headache
C0018681|T184|Cephalodynia|Headache
C0018681|T184|Headaches|Headache
C0018681|T184|ache head|Headache
C0018681|T184|cephalgias|Headache
C0018681|T184|head pain|Headache
C0018681|T184|R51|Headache
C0018681|T184|R51.9|Headache
C0231528|T184|myalgia|Muscle or body aches
C0231528|T184|myalgias|Muscle or body aches
C0231528|T184|myodynia|Muscle or body aches
C0231528|T184|Myoneuralgia|Muscle or body aches
C0231528|T184|Myosalgia|Muscle or body aches
C0231528|T184|muscle pain|Muscle or body aches
C0231528|T184|muscle pains|Muscle or body aches
C0231528|T184|muscle soreness|Muscle or body aches
C0231528|T184|aching muscles|Muscle or body aches
C0231528|T184|muscle ache|Muscle or body aches
C0231528|T184|muscle aches|Muscle or body aches
C0231528|T184|muscles aching|Muscle or body aches
C0231528|T184|aching muscles|Muscle or body aches
C0231528|T184|M79.1|Muscle or body aches
C0281856|T184|generalized aches and pains|Muscle or body aches
C0281856|T184|generalized body aches|Muscle or body aches
C0281856|T184|body aches|Muscle or body aches
C0281856|T184|aching body|Muscle or body aches
C0281856|T184|generalized pain|Muscle or body aches
C0281856|T184|generalized ache|Muscle or body aches
C0281856|T184|generalized aches|Muscle or body aches
C0281856|T184|generalized aching|Muscle or body aches
C0281856|T184|generalized body pain|Muscle or body aches
C0281856|T184|pain generalized|Muscle or body aches
C0281856|T184|body pain|Muscle or body aches
C0027497|T184|Nausea|Nausea or vomiting
C0027497|T184|nauseated|Nausea or vomiting
C0027497|T184|nauseating|Nausea or vomiting
C0027497|T184|nauseous|Nausea or vomiting
C0027497|T184|queasy|Nausea or vomiting
C0027497|T184|R11.0|Nausea or vomiting
C0042963|T184|Vomiting|Nausea or vomiting
C0042963|T184|vomit|Nausea or vomiting
C0042963|T184|vomited|Nausea or vomiting
C0042963|T184|throwing up|Nausea or vomiting
C0042963|T184|throw up|Nausea or vomiting
C0042963|T184|threw up|Nausea or vomiting
C0042963|T184|regurgitated|Nausea or vomiting
C0042963|T184|R11|Nausea or vomiting
C0042963|T184|R11.1|Nausea or vomiting
C0042963|T184|R11.10|Nausea or vomiting
C0027498|T184|Nausea and vomiting|Nausea or vomiting
C0003126|T033|Anosmia|Loss of taste or smell
C0003126|T033|Loss of smell|Loss of taste or smell
C0003126|T033|Loss of sense of smell|Loss of taste or smell
C0003126|T033|Lost sense of smell|Loss of taste or smell
C0003126|T033|Lost the sense of smell|Loss of taste or smell
C0003126|T033|Lost smell|Loss of taste or smell
C0003126|T033|No sense of smell|Loss of taste or smell
C0003126|T033|could not smell|Loss of taste or smell
C0003126|T033|R43|Loss of taste or smell
C0003126|T033|R43.0|Loss of taste or smell
C0003126|T033|Loss of smell|Loss of taste or smell
C0003126|T033|Loss of the sense of smell|Loss of taste or smell
C1332239|T184|Alterations in Smell or Taste|Loss of taste or smell
C1332239|T184|Loss of taste|Loss of taste or smell
C1332239|T184|Loss of the sense of taste|Loss of taste or smell
C1332239|T184|Lost the sense of taste|Loss of taste or smell
C1332239|T184|Lost sense of taste|Loss of taste or smell
C1332239|T184|Lost taste|Loss of taste or smell
C1332239|T184|Taste lost|Loss of taste or smell
C0013404|T184|Dyspnea|Dyspnea
C0013404|T184|difficult breathing|Dyspnea
C0013404|T184|difficulty breathing|Dyspnea
C0013404|T184|difficulty with breathing|Dyspnea
C0013404|T184|breathing difficulty|Dyspnea
C0013404|T184|breathlessness|Dyspnea
C0013404|T184|SOB|Dyspnea
C0013404|T184|shortness of breath|Dyspnea
C0013404|T184|short of breath|Dyspnea
C0013404|T184|R06|Dyspnea
C0013404|T184|R06.0|Dyspnea
C0242429|T184|Sore throat|Sore throat
C0242429|T184|throat pain|Sore throat
C0242429|T184|painful throat|Sore throat
C0242429|T184|pain in throat|Sore throat
C0242429|T184|pain in the throat|Sore throat
C0242429|T184|Pain in the pharynx|Sore throat
C0242429|T184|Pharyngeal pain|Sore throat
C0242429|T184|Throat discomfort|Sore throat
C0242429|T184|Throat soreness|Sore throat
C0242429|T184|Throat soreness|Sore throat
C0242429|T184|Pharyngitis|Sore throat
C0242429|T184|dynophagia|Sore throat
C0242429|T184|R07.0|Sore throat
